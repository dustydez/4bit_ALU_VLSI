magic
tech scmos
timestamp 1761150319
<< ab >>
rect 6 6 36 76
rect 37 75 114 76
rect 121 75 227 76
rect 233 75 310 76
rect 37 7 269 75
rect 270 7 310 75
rect 1 4 33 6
rect -63 -70 0 2
rect 2 -70 44 2
rect 46 -70 155 2
<< nwell >>
rect -4 76 38 81
rect -4 37 312 76
rect -63 -71 312 -30
<< pwell >>
rect -63 10 -24 37
rect -4 10 312 37
rect -63 -30 312 10
<< poly >>
rect 18 70 20 74
rect 25 70 27 74
rect 251 71 253 75
rect 258 71 260 75
rect 56 63 58 68
rect 63 63 65 68
rect 73 63 75 68
rect 80 63 82 68
rect 90 63 92 68
rect 110 63 112 68
rect 120 63 122 68
rect 127 63 129 68
rect 137 63 139 68
rect 144 63 146 68
rect 174 63 176 68
rect 184 63 186 68
rect 191 63 193 68
rect 201 63 203 68
rect 208 63 210 68
rect 39 56 45 58
rect 39 54 41 56
rect 43 54 45 56
rect 39 52 48 54
rect 18 47 20 50
rect 15 45 21 47
rect 15 43 17 45
rect 19 43 21 45
rect 15 41 21 43
rect 16 29 18 41
rect 25 38 27 50
rect 46 49 48 52
rect 157 56 163 58
rect 157 54 159 56
rect 161 54 163 56
rect 25 36 31 38
rect 25 34 27 36
rect 29 34 31 36
rect 25 32 31 34
rect 26 29 28 32
rect 46 23 48 43
rect 56 40 58 51
rect 63 48 65 51
rect 62 46 68 48
rect 62 44 64 46
rect 66 44 68 46
rect 62 42 68 44
rect 52 38 58 40
rect 73 38 75 51
rect 80 42 82 51
rect 52 36 54 38
rect 56 36 58 38
rect 52 34 58 36
rect 56 23 58 34
rect 63 36 75 38
rect 79 40 85 42
rect 79 38 81 40
rect 83 38 85 40
rect 79 36 85 38
rect 63 23 65 36
rect 69 30 75 32
rect 69 28 71 30
rect 73 28 75 30
rect 69 26 75 28
rect 73 23 75 26
rect 80 23 82 36
rect 90 32 92 51
rect 110 32 112 51
rect 120 42 122 51
rect 117 40 123 42
rect 117 38 119 40
rect 121 38 123 40
rect 117 36 123 38
rect 127 38 129 51
rect 137 48 139 51
rect 134 46 140 48
rect 134 44 136 46
rect 138 44 140 46
rect 134 42 140 44
rect 144 40 146 51
rect 154 52 163 54
rect 154 49 156 52
rect 238 62 240 66
rect 221 56 227 58
rect 221 54 223 56
rect 225 54 227 56
rect 144 38 150 40
rect 127 36 139 38
rect 87 30 93 32
rect 87 28 89 30
rect 91 28 93 30
rect 87 26 93 28
rect 109 30 115 32
rect 109 28 111 30
rect 113 28 115 30
rect 109 26 115 28
rect 90 23 92 26
rect 110 23 112 26
rect 120 23 122 36
rect 127 30 133 32
rect 127 28 129 30
rect 131 28 133 30
rect 127 26 133 28
rect 127 23 129 26
rect 137 23 139 36
rect 144 36 146 38
rect 148 36 150 38
rect 144 34 150 36
rect 144 23 146 34
rect 154 23 156 43
rect 174 32 176 51
rect 184 42 186 51
rect 181 40 187 42
rect 181 38 183 40
rect 185 38 187 40
rect 181 36 187 38
rect 191 38 193 51
rect 201 48 203 51
rect 198 46 204 48
rect 198 44 200 46
rect 202 44 204 46
rect 198 42 204 44
rect 208 40 210 51
rect 218 52 227 54
rect 218 49 220 52
rect 289 62 295 64
rect 289 60 291 62
rect 293 60 295 62
rect 279 55 281 60
rect 289 58 295 60
rect 208 38 214 40
rect 191 36 203 38
rect 173 30 179 32
rect 173 28 175 30
rect 177 28 179 30
rect 173 26 179 28
rect 174 23 176 26
rect 184 23 186 36
rect 191 30 197 32
rect 191 28 193 30
rect 195 28 197 30
rect 191 26 197 28
rect 191 23 193 26
rect 201 23 203 36
rect 208 36 210 38
rect 212 36 214 38
rect 208 34 214 36
rect 208 23 210 34
rect 218 23 220 43
rect 238 41 240 50
rect 251 48 253 53
rect 248 46 254 48
rect 248 44 250 46
rect 252 44 254 46
rect 248 42 254 44
rect 238 39 244 41
rect 238 37 240 39
rect 242 37 244 39
rect 238 35 244 37
rect 238 26 240 35
rect 248 26 250 42
rect 258 40 260 53
rect 289 53 291 58
rect 299 53 301 58
rect 279 40 281 43
rect 289 40 291 43
rect 258 38 264 40
rect 258 36 260 38
rect 262 36 264 38
rect 258 34 264 36
rect 279 38 285 40
rect 279 36 281 38
rect 283 36 285 38
rect 289 37 293 40
rect 279 34 285 36
rect 258 26 260 34
rect 279 26 281 34
rect 16 18 18 23
rect 26 18 28 23
rect 291 23 293 37
rect 299 32 301 43
rect 298 30 304 32
rect 298 28 300 30
rect 302 28 304 30
rect 298 26 304 28
rect 298 23 300 26
rect 46 9 48 17
rect 56 13 58 17
rect 63 9 65 17
rect 73 12 75 17
rect 80 12 82 17
rect 90 12 92 17
rect 110 12 112 17
rect 120 12 122 17
rect 127 12 129 17
rect 46 7 65 9
rect 137 9 139 17
rect 144 13 146 17
rect 154 9 156 17
rect 174 12 176 17
rect 184 12 186 17
rect 191 12 193 17
rect 137 7 156 9
rect 201 9 203 17
rect 208 13 210 17
rect 218 9 220 17
rect 238 16 240 20
rect 248 16 250 20
rect 258 16 260 20
rect 279 16 281 20
rect 201 7 220 9
rect 291 9 293 14
rect 298 9 300 14
rect -55 -2 -36 0
rect -55 -10 -53 -2
rect -45 -10 -43 -6
rect -38 -10 -36 -2
rect 54 -4 56 0
rect 65 -4 67 0
rect 72 -4 74 0
rect -28 -10 -26 -5
rect -21 -10 -19 -5
rect -11 -10 -9 -5
rect 13 -15 15 -10
rect -55 -36 -53 -16
rect -45 -27 -43 -16
rect -49 -29 -43 -27
rect -49 -31 -47 -29
rect -45 -31 -43 -29
rect -38 -29 -36 -16
rect -28 -19 -26 -16
rect -32 -21 -26 -19
rect -32 -23 -30 -21
rect -28 -23 -26 -21
rect -32 -25 -26 -23
rect -21 -29 -19 -16
rect -11 -19 -9 -16
rect -14 -21 -8 -19
rect -14 -23 -12 -21
rect -10 -23 -8 -21
rect -14 -25 -8 -23
rect 23 -18 25 -13
rect 33 -18 35 -13
rect -38 -31 -26 -29
rect -49 -33 -43 -31
rect -55 -45 -53 -42
rect -62 -47 -53 -45
rect -45 -44 -43 -33
rect -39 -37 -33 -35
rect -39 -39 -37 -37
rect -35 -39 -33 -37
rect -39 -41 -33 -39
rect -38 -44 -36 -41
rect -28 -44 -26 -31
rect -22 -31 -16 -29
rect -22 -33 -20 -31
rect -18 -33 -16 -31
rect -22 -35 -16 -33
rect -21 -44 -19 -35
rect -11 -44 -9 -25
rect 13 -27 15 -24
rect 23 -27 25 -24
rect 13 -29 19 -27
rect 13 -31 15 -29
rect 17 -31 19 -29
rect 13 -33 19 -31
rect 23 -29 29 -27
rect 23 -31 25 -29
rect 27 -31 29 -29
rect 23 -33 29 -31
rect 13 -36 15 -33
rect -62 -49 -60 -47
rect -58 -49 -56 -47
rect -62 -51 -56 -49
rect 26 -43 28 -33
rect 33 -34 35 -24
rect 54 -27 56 -18
rect 92 -10 94 -5
rect 102 -10 104 -5
rect 112 -7 114 -2
rect 122 -4 124 0
rect 143 -4 145 0
rect 154 -4 156 0
rect 161 -4 163 0
rect 65 -27 67 -24
rect 72 -27 74 -24
rect 92 -27 94 -24
rect 102 -27 104 -24
rect 52 -29 58 -27
rect 52 -31 54 -29
rect 56 -31 58 -29
rect 52 -33 58 -31
rect 62 -29 68 -27
rect 62 -31 64 -29
rect 66 -31 68 -29
rect 62 -33 68 -31
rect 72 -29 94 -27
rect 72 -31 74 -29
rect 76 -31 81 -29
rect 83 -31 94 -29
rect 72 -33 94 -31
rect 98 -29 104 -27
rect 98 -31 100 -29
rect 102 -31 104 -29
rect 98 -33 104 -31
rect 112 -30 114 -17
rect 122 -20 124 -17
rect 118 -22 124 -20
rect 118 -24 120 -22
rect 122 -24 124 -22
rect 118 -26 124 -24
rect 112 -32 118 -30
rect 33 -36 39 -34
rect 54 -36 56 -33
rect 64 -36 66 -33
rect 74 -36 76 -33
rect 92 -36 94 -33
rect 99 -36 101 -33
rect 112 -34 114 -32
rect 116 -34 118 -32
rect 109 -36 118 -34
rect 33 -38 35 -36
rect 37 -38 39 -36
rect 33 -40 39 -38
rect 33 -43 35 -40
rect -45 -61 -43 -56
rect -38 -61 -36 -56
rect -28 -61 -26 -56
rect -21 -61 -19 -56
rect -11 -61 -9 -56
rect 13 -59 15 -54
rect 109 -39 111 -36
rect 122 -39 124 -26
rect 143 -27 145 -18
rect 181 -10 183 -5
rect 191 -10 193 -5
rect 201 -7 203 -2
rect 211 -4 213 0
rect 231 -2 250 0
rect 231 -12 233 -2
rect 241 -10 243 -6
rect 248 -10 250 -2
rect 258 -10 260 -5
rect 265 -10 267 -5
rect 275 -10 277 -5
rect 154 -27 156 -24
rect 161 -27 163 -24
rect 181 -27 183 -24
rect 191 -27 193 -24
rect 141 -29 147 -27
rect 141 -31 143 -29
rect 145 -31 147 -29
rect 141 -33 147 -31
rect 151 -29 157 -27
rect 151 -31 153 -29
rect 155 -31 157 -29
rect 151 -33 157 -31
rect 161 -29 183 -27
rect 161 -31 163 -29
rect 165 -31 170 -29
rect 172 -31 183 -29
rect 161 -33 183 -31
rect 187 -29 193 -27
rect 187 -31 189 -29
rect 191 -31 193 -29
rect 187 -33 193 -31
rect 201 -30 203 -17
rect 211 -20 213 -17
rect 207 -22 213 -20
rect 207 -24 209 -22
rect 211 -24 213 -22
rect 207 -26 213 -24
rect 201 -32 207 -30
rect 143 -36 145 -33
rect 153 -36 155 -33
rect 163 -36 165 -33
rect 181 -36 183 -33
rect 188 -36 190 -33
rect 201 -34 203 -32
rect 205 -34 207 -32
rect 198 -36 207 -34
rect 109 -57 111 -52
rect 26 -68 28 -64
rect 33 -68 35 -64
rect 54 -68 56 -64
rect 64 -68 66 -64
rect 74 -68 76 -64
rect 92 -66 94 -61
rect 99 -66 101 -61
rect 198 -39 200 -36
rect 211 -39 213 -26
rect 231 -36 233 -18
rect 241 -27 243 -18
rect 237 -29 243 -27
rect 237 -31 239 -29
rect 241 -31 243 -29
rect 237 -33 243 -31
rect 248 -31 250 -18
rect 258 -21 260 -18
rect 254 -23 260 -21
rect 254 -25 256 -23
rect 258 -25 260 -23
rect 254 -27 260 -25
rect 248 -33 260 -31
rect 265 -32 267 -18
rect 295 -15 297 -10
rect 275 -22 277 -19
rect 272 -24 278 -22
rect 272 -26 274 -24
rect 276 -26 278 -24
rect 272 -28 278 -26
rect 295 -27 297 -24
rect 198 -57 200 -52
rect 122 -68 124 -64
rect 143 -68 145 -64
rect 153 -68 155 -64
rect 163 -68 165 -64
rect 181 -66 183 -61
rect 188 -66 190 -61
rect 231 -47 233 -44
rect 224 -49 233 -47
rect 241 -48 243 -33
rect 247 -39 253 -37
rect 247 -41 249 -39
rect 251 -41 253 -39
rect 247 -43 253 -41
rect 248 -48 250 -43
rect 258 -48 260 -33
rect 264 -34 270 -32
rect 264 -36 266 -34
rect 268 -36 270 -34
rect 264 -38 270 -36
rect 265 -48 267 -38
rect 275 -46 277 -28
rect 295 -29 301 -27
rect 295 -31 297 -29
rect 299 -31 301 -29
rect 295 -33 301 -31
rect 295 -36 297 -33
rect 224 -51 226 -49
rect 228 -51 230 -49
rect 224 -53 230 -51
rect 295 -59 297 -54
rect 211 -68 213 -64
rect 241 -68 243 -64
rect 248 -68 250 -64
rect 258 -68 260 -64
rect 265 -68 267 -64
rect 275 -68 277 -64
<< ndif >>
rect 8 27 16 29
rect 8 25 10 27
rect 12 25 16 27
rect 8 23 16 25
rect 18 27 26 29
rect 18 25 21 27
rect 23 25 26 27
rect 18 23 26 25
rect 28 27 35 29
rect 28 25 31 27
rect 33 25 35 27
rect 28 23 35 25
rect 231 24 238 26
rect 39 21 46 23
rect 39 19 41 21
rect 43 19 46 21
rect 39 17 46 19
rect 48 21 56 23
rect 48 19 51 21
rect 53 19 56 21
rect 48 17 56 19
rect 58 17 63 23
rect 65 21 73 23
rect 65 19 68 21
rect 70 19 73 21
rect 65 17 73 19
rect 75 17 80 23
rect 82 21 90 23
rect 82 19 85 21
rect 87 19 90 21
rect 82 17 90 19
rect 92 21 99 23
rect 92 19 95 21
rect 97 19 99 21
rect 92 17 99 19
rect 103 21 110 23
rect 103 19 105 21
rect 107 19 110 21
rect 103 17 110 19
rect 112 21 120 23
rect 112 19 115 21
rect 117 19 120 21
rect 112 17 120 19
rect 122 17 127 23
rect 129 21 137 23
rect 129 19 132 21
rect 134 19 137 21
rect 129 17 137 19
rect 139 17 144 23
rect 146 21 154 23
rect 146 19 149 21
rect 151 19 154 21
rect 146 17 154 19
rect 156 21 163 23
rect 156 19 159 21
rect 161 19 163 21
rect 156 17 163 19
rect 167 21 174 23
rect 167 19 169 21
rect 171 19 174 21
rect 167 17 174 19
rect 176 21 184 23
rect 176 19 179 21
rect 181 19 184 21
rect 176 17 184 19
rect 186 17 191 23
rect 193 21 201 23
rect 193 19 196 21
rect 198 19 201 21
rect 193 17 201 19
rect 203 17 208 23
rect 210 21 218 23
rect 210 19 213 21
rect 215 19 218 21
rect 210 17 218 19
rect 220 21 227 23
rect 220 19 223 21
rect 225 19 227 21
rect 231 22 233 24
rect 235 22 238 24
rect 231 20 238 22
rect 240 24 248 26
rect 240 22 243 24
rect 245 22 248 24
rect 240 20 248 22
rect 250 24 258 26
rect 250 22 253 24
rect 255 22 258 24
rect 250 20 258 22
rect 260 24 267 26
rect 260 22 263 24
rect 265 22 267 24
rect 260 20 267 22
rect 272 24 279 26
rect 272 22 274 24
rect 276 22 279 24
rect 272 20 279 22
rect 281 23 289 26
rect 281 20 291 23
rect 220 17 227 19
rect 283 14 291 20
rect 293 14 298 23
rect 300 21 307 23
rect 300 19 303 21
rect 305 19 307 21
rect 300 17 307 19
rect 300 14 305 17
rect 283 12 289 14
rect 283 10 285 12
rect 287 10 289 12
rect 283 8 289 10
rect 17 -7 23 -5
rect 17 -9 19 -7
rect 21 -9 23 -7
rect -62 -12 -55 -10
rect -62 -14 -60 -12
rect -58 -14 -55 -12
rect -62 -16 -55 -14
rect -53 -12 -45 -10
rect -53 -14 -50 -12
rect -48 -14 -45 -12
rect -53 -16 -45 -14
rect -43 -16 -38 -10
rect -36 -12 -28 -10
rect -36 -14 -33 -12
rect -31 -14 -28 -12
rect -36 -16 -28 -14
rect -26 -16 -21 -10
rect -19 -12 -11 -10
rect -19 -14 -16 -12
rect -14 -14 -11 -12
rect -19 -16 -11 -14
rect -9 -12 -2 -10
rect -9 -14 -6 -12
rect -4 -14 -2 -12
rect -9 -16 -2 -14
rect 17 -11 23 -9
rect 36 -7 42 -5
rect 36 -9 38 -7
rect 40 -9 42 -7
rect 36 -11 42 -9
rect 49 -11 54 -4
rect 17 -15 21 -11
rect 8 -18 13 -15
rect 6 -20 13 -18
rect 6 -22 8 -20
rect 10 -22 13 -20
rect 6 -24 13 -22
rect 15 -18 21 -15
rect 37 -18 42 -11
rect 47 -13 54 -11
rect 47 -15 49 -13
rect 51 -15 54 -13
rect 47 -18 54 -15
rect 56 -6 65 -4
rect 56 -8 60 -6
rect 62 -8 65 -6
rect 56 -18 65 -8
rect 15 -24 23 -18
rect 25 -20 33 -18
rect 25 -22 28 -20
rect 30 -22 33 -20
rect 25 -24 33 -22
rect 35 -24 42 -18
rect 58 -24 65 -18
rect 67 -24 72 -4
rect 74 -11 79 -4
rect 117 -7 122 -4
rect 107 -10 112 -7
rect 74 -13 81 -11
rect 74 -15 77 -13
rect 79 -15 81 -13
rect 74 -17 81 -15
rect 85 -13 92 -10
rect 85 -15 87 -13
rect 89 -15 92 -13
rect 74 -24 79 -17
rect 85 -20 92 -15
rect 85 -22 87 -20
rect 89 -22 92 -20
rect 85 -24 92 -22
rect 94 -20 102 -10
rect 94 -22 97 -20
rect 99 -22 102 -20
rect 94 -24 102 -22
rect 104 -12 112 -10
rect 104 -14 107 -12
rect 109 -14 112 -12
rect 104 -17 112 -14
rect 114 -9 122 -7
rect 114 -11 117 -9
rect 119 -11 122 -9
rect 114 -17 122 -11
rect 124 -11 129 -4
rect 138 -11 143 -4
rect 124 -13 131 -11
rect 124 -15 127 -13
rect 129 -15 131 -13
rect 124 -17 131 -15
rect 136 -13 143 -11
rect 136 -15 138 -13
rect 140 -15 143 -13
rect 104 -24 109 -17
rect 136 -18 143 -15
rect 145 -6 154 -4
rect 145 -8 149 -6
rect 151 -8 154 -6
rect 145 -18 154 -8
rect 147 -24 154 -18
rect 156 -24 161 -4
rect 163 -11 168 -4
rect 206 -7 211 -4
rect 196 -10 201 -7
rect 163 -13 170 -11
rect 163 -15 166 -13
rect 168 -15 170 -13
rect 163 -17 170 -15
rect 174 -13 181 -10
rect 174 -15 176 -13
rect 178 -15 181 -13
rect 163 -24 168 -17
rect 174 -20 181 -15
rect 174 -22 176 -20
rect 178 -22 181 -20
rect 174 -24 181 -22
rect 183 -20 191 -10
rect 183 -22 186 -20
rect 188 -22 191 -20
rect 183 -24 191 -22
rect 193 -12 201 -10
rect 193 -14 196 -12
rect 198 -14 201 -12
rect 193 -17 201 -14
rect 203 -9 211 -7
rect 203 -11 206 -9
rect 208 -11 211 -9
rect 203 -17 211 -11
rect 213 -11 218 -4
rect 213 -13 220 -11
rect 235 -12 241 -10
rect 213 -15 216 -13
rect 218 -15 220 -13
rect 213 -17 220 -15
rect 224 -14 231 -12
rect 224 -16 226 -14
rect 228 -16 231 -14
rect 193 -24 198 -17
rect 224 -18 231 -16
rect 233 -14 241 -12
rect 233 -16 236 -14
rect 238 -16 241 -14
rect 233 -18 241 -16
rect 243 -18 248 -10
rect 250 -12 258 -10
rect 250 -14 253 -12
rect 255 -14 258 -12
rect 250 -18 258 -14
rect 260 -18 265 -10
rect 267 -12 275 -10
rect 267 -14 270 -12
rect 272 -14 275 -12
rect 267 -18 275 -14
rect 270 -19 275 -18
rect 277 -13 282 -10
rect 277 -15 284 -13
rect 277 -17 280 -15
rect 282 -17 284 -15
rect 277 -19 284 -17
rect 290 -18 295 -15
rect 288 -20 295 -18
rect 288 -22 290 -20
rect 292 -22 295 -20
rect 288 -24 295 -22
rect 297 -17 308 -15
rect 297 -19 304 -17
rect 306 -19 308 -17
rect 297 -24 308 -19
<< pdif >>
rect 13 64 18 70
rect 11 62 18 64
rect 11 60 13 62
rect 15 60 18 62
rect 11 58 18 60
rect 13 50 18 58
rect 20 50 25 70
rect 27 68 36 70
rect 242 69 251 71
rect 27 66 32 68
rect 34 66 36 68
rect 27 61 36 66
rect 242 67 245 69
rect 247 67 251 69
rect 27 59 32 61
rect 34 59 36 61
rect 27 56 36 59
rect 49 61 56 63
rect 49 59 51 61
rect 53 59 56 61
rect 49 57 56 59
rect 27 50 35 56
rect 50 51 56 57
rect 58 51 63 63
rect 65 55 73 63
rect 65 53 68 55
rect 70 53 73 55
rect 65 51 73 53
rect 75 51 80 63
rect 82 61 90 63
rect 82 59 85 61
rect 87 59 90 61
rect 82 51 90 59
rect 92 57 97 63
rect 105 57 110 63
rect 92 55 99 57
rect 92 53 95 55
rect 97 53 99 55
rect 92 51 99 53
rect 103 55 110 57
rect 103 53 105 55
rect 107 53 110 55
rect 103 51 110 53
rect 112 61 120 63
rect 112 59 115 61
rect 117 59 120 61
rect 112 51 120 59
rect 122 51 127 63
rect 129 55 137 63
rect 129 53 132 55
rect 134 53 137 55
rect 129 51 137 53
rect 139 51 144 63
rect 146 61 153 63
rect 146 59 149 61
rect 151 59 153 61
rect 146 57 153 59
rect 146 51 152 57
rect 169 57 174 63
rect 50 49 54 51
rect 39 47 46 49
rect 39 45 41 47
rect 43 45 46 47
rect 39 43 46 45
rect 48 43 54 49
rect 148 49 152 51
rect 167 55 174 57
rect 167 53 169 55
rect 171 53 174 55
rect 167 51 174 53
rect 176 61 184 63
rect 176 59 179 61
rect 181 59 184 61
rect 176 51 184 59
rect 186 51 191 63
rect 193 55 201 63
rect 193 53 196 55
rect 198 53 201 55
rect 193 51 201 53
rect 203 51 208 63
rect 210 61 217 63
rect 242 62 251 67
rect 210 59 213 61
rect 215 59 217 61
rect 210 57 217 59
rect 231 60 238 62
rect 231 58 233 60
rect 235 58 238 60
rect 210 51 216 57
rect 231 56 238 58
rect 148 43 154 49
rect 156 47 163 49
rect 156 45 159 47
rect 161 45 163 47
rect 156 43 163 45
rect 212 49 216 51
rect 233 50 238 56
rect 240 53 251 62
rect 253 53 258 71
rect 260 64 265 71
rect 260 62 267 64
rect 260 60 263 62
rect 265 60 267 62
rect 260 58 267 60
rect 260 53 265 58
rect 240 50 248 53
rect 212 43 218 49
rect 220 47 227 49
rect 220 45 223 47
rect 225 45 227 47
rect 220 43 227 45
rect 274 49 279 55
rect 272 47 279 49
rect 272 45 274 47
rect 276 45 279 47
rect 272 43 279 45
rect 281 53 287 55
rect 281 47 289 53
rect 281 45 284 47
rect 286 45 289 47
rect 281 43 289 45
rect 291 47 299 53
rect 291 45 294 47
rect 296 45 299 47
rect 291 43 299 45
rect 301 51 308 53
rect 301 49 304 51
rect 306 49 308 51
rect 301 43 308 49
rect -62 -38 -55 -36
rect -62 -40 -60 -38
rect -58 -40 -55 -38
rect -62 -42 -55 -40
rect -53 -42 -47 -36
rect -51 -44 -47 -42
rect 8 -41 13 -36
rect 6 -43 13 -41
rect -51 -50 -45 -44
rect -52 -52 -45 -50
rect -52 -54 -50 -52
rect -48 -54 -45 -52
rect -52 -56 -45 -54
rect -43 -56 -38 -44
rect -36 -46 -28 -44
rect -36 -48 -33 -46
rect -31 -48 -28 -46
rect -36 -56 -28 -48
rect -26 -56 -21 -44
rect -19 -52 -11 -44
rect -19 -54 -16 -52
rect -14 -54 -11 -52
rect -19 -56 -11 -54
rect -9 -46 -2 -44
rect -9 -48 -6 -46
rect -4 -48 -2 -46
rect -9 -50 -2 -48
rect 6 -45 8 -43
rect 10 -45 13 -43
rect 6 -50 13 -45
rect -9 -56 -4 -50
rect 6 -52 8 -50
rect 10 -52 13 -50
rect 6 -54 13 -52
rect 15 -43 23 -36
rect 47 -38 54 -36
rect 47 -40 49 -38
rect 51 -40 54 -38
rect 15 -54 26 -43
rect 17 -60 26 -54
rect 17 -62 19 -60
rect 21 -62 26 -60
rect 17 -64 26 -62
rect 28 -64 33 -43
rect 35 -51 40 -43
rect 47 -45 54 -40
rect 47 -47 49 -45
rect 51 -47 54 -45
rect 47 -49 54 -47
rect 35 -53 42 -51
rect 35 -55 38 -53
rect 40 -55 42 -53
rect 35 -57 42 -55
rect 35 -64 40 -57
rect 49 -64 54 -49
rect 56 -53 64 -36
rect 56 -55 59 -53
rect 61 -55 64 -53
rect 56 -60 64 -55
rect 56 -62 59 -60
rect 61 -62 64 -60
rect 56 -64 64 -62
rect 66 -45 74 -36
rect 66 -47 69 -45
rect 71 -47 74 -45
rect 66 -52 74 -47
rect 66 -54 69 -52
rect 71 -54 74 -52
rect 66 -64 74 -54
rect 76 -53 92 -36
rect 76 -55 81 -53
rect 83 -55 92 -53
rect 76 -60 92 -55
rect 76 -62 81 -60
rect 83 -61 92 -60
rect 94 -61 99 -36
rect 101 -39 106 -36
rect 136 -38 143 -36
rect 101 -41 109 -39
rect 101 -43 104 -41
rect 106 -43 109 -41
rect 101 -52 109 -43
rect 111 -52 122 -39
rect 101 -61 106 -52
rect 113 -60 122 -52
rect 83 -62 90 -61
rect 76 -64 90 -62
rect 113 -62 116 -60
rect 118 -62 122 -60
rect 113 -64 122 -62
rect 124 -41 131 -39
rect 124 -43 127 -41
rect 129 -43 131 -41
rect 124 -48 131 -43
rect 124 -50 127 -48
rect 129 -50 131 -48
rect 136 -40 138 -38
rect 140 -40 143 -38
rect 136 -45 143 -40
rect 136 -47 138 -45
rect 140 -47 143 -45
rect 136 -49 143 -47
rect 124 -52 131 -50
rect 124 -64 129 -52
rect 138 -64 143 -49
rect 145 -53 153 -36
rect 145 -55 148 -53
rect 150 -55 153 -53
rect 145 -60 153 -55
rect 145 -62 148 -60
rect 150 -62 153 -60
rect 145 -64 153 -62
rect 155 -45 163 -36
rect 155 -47 158 -45
rect 160 -47 163 -45
rect 155 -52 163 -47
rect 155 -54 158 -52
rect 160 -54 163 -52
rect 155 -64 163 -54
rect 165 -53 181 -36
rect 165 -55 170 -53
rect 172 -55 181 -53
rect 165 -60 181 -55
rect 165 -62 170 -60
rect 172 -61 181 -60
rect 183 -61 188 -36
rect 190 -39 195 -36
rect 224 -38 231 -36
rect 190 -41 198 -39
rect 190 -43 193 -41
rect 195 -43 198 -41
rect 190 -52 198 -43
rect 200 -52 211 -39
rect 190 -61 195 -52
rect 202 -60 211 -52
rect 172 -62 179 -61
rect 165 -64 179 -62
rect 202 -62 205 -60
rect 207 -62 211 -60
rect 202 -64 211 -62
rect 213 -41 220 -39
rect 213 -43 216 -41
rect 218 -43 220 -41
rect 224 -40 226 -38
rect 228 -40 231 -38
rect 224 -42 231 -40
rect 213 -48 220 -43
rect 226 -44 231 -42
rect 233 -44 239 -36
rect 213 -50 216 -48
rect 218 -50 220 -48
rect 213 -52 220 -50
rect 235 -48 239 -44
rect 288 -38 295 -36
rect 288 -40 290 -38
rect 292 -40 295 -38
rect 288 -45 295 -40
rect 270 -48 275 -46
rect 213 -64 218 -52
rect 235 -52 241 -48
rect 234 -60 241 -52
rect 234 -62 236 -60
rect 238 -62 241 -60
rect 234 -64 241 -62
rect 243 -64 248 -48
rect 250 -50 258 -48
rect 250 -52 253 -50
rect 255 -52 258 -50
rect 250 -64 258 -52
rect 260 -64 265 -48
rect 267 -60 275 -48
rect 267 -62 270 -60
rect 272 -62 275 -60
rect 267 -64 275 -62
rect 277 -51 282 -46
rect 288 -47 290 -45
rect 292 -47 295 -45
rect 288 -49 295 -47
rect 277 -53 284 -51
rect 277 -55 280 -53
rect 282 -55 284 -53
rect 290 -54 295 -49
rect 297 -53 306 -36
rect 297 -54 301 -53
rect 277 -57 284 -55
rect 277 -64 282 -57
rect 299 -55 301 -54
rect 303 -55 306 -53
rect 299 -57 306 -55
<< alu1 >>
rect 5 72 327 76
rect 5 70 42 72
rect 44 70 158 72
rect 160 70 222 72
rect 224 70 234 72
rect 236 70 275 72
rect 277 70 289 72
rect 291 70 303 72
rect 305 70 327 72
rect 5 69 327 70
rect 5 68 36 69
rect 8 62 17 63
rect 8 60 13 62
rect 15 60 17 62
rect 8 59 17 60
rect 8 42 12 59
rect 39 61 44 63
rect 39 59 40 61
rect 42 59 44 61
rect 39 56 44 59
rect 158 60 163 64
rect 158 58 160 60
rect 162 58 163 60
rect 227 68 231 69
rect 222 61 227 64
rect 222 59 224 61
rect 226 59 227 61
rect 158 56 163 58
rect 222 56 227 59
rect 24 54 28 55
rect 24 52 25 54
rect 27 52 28 54
rect 24 50 28 52
rect 39 54 41 56
rect 43 55 44 56
rect 93 55 99 56
rect 43 54 52 55
rect 39 51 52 54
rect 86 53 95 55
rect 97 53 99 55
rect 86 51 99 53
rect 8 40 9 42
rect 11 40 12 42
rect 16 46 28 50
rect 32 46 36 47
rect 16 45 20 46
rect 16 43 17 45
rect 19 43 20 45
rect 16 41 20 43
rect 32 44 33 46
rect 35 44 36 46
rect 8 37 12 40
rect 32 39 36 44
rect 8 33 20 37
rect 24 36 36 39
rect 24 34 27 36
rect 29 34 36 36
rect 24 33 36 34
rect 16 28 20 33
rect 16 27 25 28
rect 16 25 21 27
rect 23 25 25 27
rect 16 24 25 25
rect 53 38 59 40
rect 53 36 54 38
rect 56 36 59 38
rect 53 32 59 36
rect 47 30 59 32
rect 47 28 53 30
rect 55 28 59 30
rect 47 26 59 28
rect 70 41 76 47
rect 70 40 85 41
rect 70 39 81 40
rect 70 37 76 39
rect 78 38 81 39
rect 83 38 85 40
rect 78 37 85 38
rect 70 35 85 37
rect 95 39 99 51
rect 95 37 96 39
rect 98 37 99 39
rect 95 22 99 37
rect 93 21 99 22
rect 93 19 95 21
rect 97 19 99 21
rect 93 18 99 19
rect 103 55 109 56
rect 158 55 159 56
rect 103 53 105 55
rect 107 53 116 55
rect 103 51 116 53
rect 150 54 159 55
rect 161 54 163 56
rect 150 51 163 54
rect 167 55 173 56
rect 222 55 223 56
rect 167 53 169 55
rect 171 53 180 55
rect 167 51 180 53
rect 214 54 223 55
rect 225 54 227 56
rect 214 51 227 54
rect 231 60 244 63
rect 231 58 233 60
rect 235 59 244 60
rect 103 22 107 51
rect 126 41 132 47
rect 117 40 132 41
rect 117 38 119 40
rect 121 39 132 40
rect 121 38 124 39
rect 117 37 124 38
rect 126 37 132 39
rect 117 35 132 37
rect 143 38 149 40
rect 143 36 146 38
rect 148 36 149 38
rect 143 32 149 36
rect 143 30 155 32
rect 143 28 148 30
rect 150 28 155 30
rect 143 26 155 28
rect 103 21 109 22
rect 103 19 105 21
rect 107 19 109 21
rect 103 18 109 19
rect 167 30 171 51
rect 167 28 168 30
rect 170 28 171 30
rect 167 22 171 28
rect 190 42 196 47
rect 190 41 193 42
rect 181 40 193 41
rect 195 40 196 42
rect 181 38 183 40
rect 185 38 196 40
rect 181 35 196 38
rect 207 38 213 40
rect 207 36 210 38
rect 212 36 213 38
rect 207 32 213 36
rect 207 29 219 32
rect 207 27 216 29
rect 218 27 219 29
rect 207 26 219 27
rect 167 21 173 22
rect 167 19 169 21
rect 171 19 173 21
rect 167 18 173 19
rect 231 42 235 58
rect 231 40 232 42
rect 234 40 235 42
rect 231 26 235 40
rect 255 55 259 56
rect 255 53 256 55
rect 258 53 259 55
rect 255 47 259 53
rect 246 46 259 47
rect 246 44 250 46
rect 252 44 259 46
rect 246 43 259 44
rect 263 39 267 48
rect 254 38 267 39
rect 254 36 260 38
rect 262 36 264 38
rect 266 36 267 38
rect 254 35 267 36
rect 263 34 267 35
rect 272 47 276 56
rect 272 45 274 47
rect 231 24 236 26
rect 231 22 233 24
rect 235 22 236 24
rect 231 18 236 22
rect 272 29 276 45
rect 287 62 300 64
rect 287 60 291 62
rect 293 60 300 62
rect 287 58 300 60
rect 287 55 293 58
rect 287 53 289 55
rect 291 53 293 55
rect 287 51 293 53
rect 304 38 308 40
rect 304 36 305 38
rect 307 36 308 38
rect 272 27 273 29
rect 275 27 276 29
rect 272 24 276 27
rect 272 22 274 24
rect 276 22 284 24
rect 272 18 284 22
rect 304 31 308 36
rect 295 30 308 31
rect 295 28 300 30
rect 302 28 308 30
rect 295 26 308 28
rect 0 12 312 13
rect -1 11 234 12
rect -1 9 11 11
rect 13 9 31 11
rect 33 10 234 11
rect 236 10 262 12
rect 264 10 275 12
rect 277 10 285 12
rect 287 10 312 12
rect 33 9 312 10
rect -1 5 312 9
rect -63 -3 312 5
rect -63 -5 9 -3
rect 11 -5 291 -3
rect 293 -5 303 -3
rect 305 -5 312 -3
rect -63 -6 312 -5
rect -8 -12 -2 -11
rect -8 -14 -6 -12
rect -4 -14 -2 -12
rect -8 -15 -2 -14
rect -54 -20 -42 -19
rect -54 -22 -50 -20
rect -48 -22 -42 -20
rect -54 -25 -42 -22
rect -48 -29 -42 -25
rect -48 -31 -47 -29
rect -45 -31 -42 -29
rect -48 -33 -42 -31
rect -31 -31 -16 -28
rect -31 -33 -29 -31
rect -27 -33 -20 -31
rect -18 -33 -16 -31
rect -31 -34 -16 -33
rect -31 -40 -25 -34
rect -6 -44 -2 -15
rect 46 -13 68 -12
rect 46 -15 49 -13
rect 51 -15 68 -13
rect 46 -16 68 -15
rect 126 -13 131 -11
rect 126 -15 127 -13
rect 129 -15 131 -13
rect -62 -47 -49 -44
rect -62 -49 -60 -47
rect -58 -48 -49 -47
rect -15 -46 -2 -44
rect -15 -48 -6 -46
rect -4 -48 -2 -46
rect -58 -49 -57 -48
rect -8 -49 -2 -48
rect 6 -20 11 -18
rect 6 -22 8 -20
rect 10 -22 11 -20
rect 6 -24 11 -22
rect 38 -20 42 -19
rect 38 -22 39 -20
rect 41 -22 42 -20
rect 6 -31 10 -24
rect 6 -33 7 -31
rect 9 -33 10 -31
rect 6 -43 10 -33
rect 38 -28 42 -22
rect 6 -45 8 -43
rect -62 -53 -57 -49
rect 6 -50 10 -45
rect -62 -55 -60 -53
rect -58 -55 -57 -53
rect -62 -57 -57 -55
rect 6 -52 8 -50
rect 21 -29 42 -28
rect 21 -31 25 -29
rect 27 -31 42 -29
rect 21 -32 42 -31
rect 46 -36 50 -16
rect 21 -38 35 -36
rect 37 -38 42 -36
rect 21 -40 42 -38
rect 38 -42 42 -40
rect 46 -38 52 -36
rect 46 -40 49 -38
rect 51 -40 52 -38
rect 46 -42 52 -40
rect 38 -45 52 -42
rect 38 -46 49 -45
rect 38 -49 42 -46
rect 46 -47 49 -46
rect 51 -47 52 -45
rect 46 -49 52 -47
rect 79 -28 83 -19
rect 126 -17 131 -15
rect 70 -29 85 -28
rect 70 -31 74 -29
rect 76 -31 81 -29
rect 83 -31 85 -29
rect 70 -32 85 -31
rect 95 -29 103 -27
rect 95 -31 96 -29
rect 98 -31 100 -29
rect 102 -31 103 -29
rect 95 -33 103 -31
rect 95 -36 100 -33
rect 62 -40 100 -36
rect 127 -37 131 -17
rect 127 -39 128 -37
rect 130 -39 131 -37
rect 126 -41 131 -39
rect 126 -43 127 -41
rect 129 -43 131 -41
rect 126 -48 131 -43
rect 126 -50 127 -48
rect 129 -50 131 -48
rect 135 -13 157 -12
rect 135 -15 138 -13
rect 140 -15 157 -13
rect 135 -16 157 -15
rect 215 -13 220 -11
rect 215 -15 216 -13
rect 218 -15 220 -13
rect 135 -20 139 -16
rect 135 -22 136 -20
rect 138 -22 139 -20
rect 135 -36 139 -22
rect 168 -20 172 -19
rect 168 -22 169 -20
rect 171 -22 172 -20
rect 135 -38 141 -36
rect 135 -40 138 -38
rect 140 -40 141 -38
rect 135 -45 141 -40
rect 135 -47 138 -45
rect 140 -47 141 -45
rect 135 -49 141 -47
rect 168 -28 172 -22
rect 215 -17 220 -15
rect 216 -19 217 -17
rect 219 -19 220 -17
rect 159 -29 174 -28
rect 159 -31 163 -29
rect 165 -31 170 -29
rect 172 -31 174 -29
rect 159 -32 174 -31
rect 184 -29 192 -27
rect 184 -31 189 -29
rect 191 -31 192 -29
rect 184 -33 192 -31
rect 184 -36 189 -33
rect 151 -37 189 -36
rect 151 -39 158 -37
rect 160 -39 189 -37
rect 151 -40 189 -39
rect 216 -39 220 -19
rect 215 -41 220 -39
rect 280 -13 284 -11
rect 279 -15 284 -13
rect 279 -17 280 -15
rect 282 -17 284 -15
rect 279 -19 284 -17
rect 231 -21 244 -20
rect 231 -23 241 -21
rect 243 -23 244 -21
rect 231 -24 244 -23
rect 238 -29 244 -24
rect 238 -31 239 -29
rect 241 -31 244 -29
rect 238 -33 244 -31
rect 264 -34 268 -27
rect 264 -35 266 -34
rect 256 -36 266 -35
rect 256 -37 268 -36
rect 256 -39 261 -37
rect 263 -39 268 -37
rect 256 -41 268 -39
rect 215 -43 216 -41
rect 218 -43 220 -41
rect 215 -48 220 -43
rect 126 -52 131 -50
rect 215 -50 216 -48
rect 218 -50 220 -48
rect 215 -52 220 -50
rect 6 -56 19 -52
rect 6 -57 10 -56
rect 118 -56 131 -52
rect 207 -56 220 -52
rect 224 -48 237 -44
rect 224 -49 229 -48
rect 280 -29 284 -19
rect 280 -31 281 -29
rect 283 -31 284 -29
rect 224 -51 226 -49
rect 228 -51 229 -49
rect 224 -57 229 -51
rect 280 -52 284 -31
rect 288 -20 292 -11
rect 288 -22 290 -20
rect 288 -24 292 -22
rect 288 -26 289 -24
rect 291 -26 292 -24
rect 288 -38 292 -26
rect 296 -27 300 -19
rect 296 -29 308 -27
rect 296 -31 297 -29
rect 299 -31 304 -29
rect 306 -31 308 -29
rect 296 -33 308 -31
rect 288 -40 290 -38
rect 288 -43 292 -40
rect 288 -45 300 -43
rect 288 -47 290 -45
rect 292 -47 300 -45
rect 288 -49 300 -47
rect 271 -53 284 -52
rect 271 -55 280 -53
rect 282 -55 284 -53
rect 271 -56 284 -55
rect -63 -63 312 -62
rect 319 -63 327 69
rect -63 -65 -59 -63
rect -57 -65 9 -63
rect 11 -65 291 -63
rect 293 -65 303 -63
rect 305 -65 327 -63
rect -63 -70 327 -65
<< alu2 >>
rect 148 65 171 69
rect 148 62 152 65
rect 24 61 152 62
rect 167 62 171 65
rect 167 61 227 62
rect 24 59 40 61
rect 42 59 152 61
rect 24 58 152 59
rect 157 60 163 61
rect 157 58 160 60
rect 162 58 163 60
rect 167 59 224 61
rect 226 59 227 61
rect 167 58 227 59
rect 24 54 28 58
rect 157 54 163 58
rect 24 52 25 54
rect 27 52 28 54
rect 24 51 28 52
rect 32 50 163 54
rect 254 55 293 56
rect 254 53 256 55
rect 258 53 289 55
rect 291 53 293 55
rect 254 52 293 53
rect 32 46 36 50
rect 254 47 259 52
rect 8 42 12 45
rect 32 44 33 46
rect 35 44 36 46
rect 32 42 36 44
rect 246 46 259 47
rect 246 44 247 46
rect 249 44 259 46
rect 246 43 259 44
rect 191 42 235 43
rect 8 40 9 42
rect 11 40 12 42
rect 8 5 12 40
rect 73 39 85 41
rect 73 37 76 39
rect 78 37 85 39
rect 73 35 85 37
rect 95 39 132 41
rect 191 40 193 42
rect 195 40 232 42
rect 234 40 235 42
rect 191 39 235 40
rect 95 37 96 39
rect 98 37 124 39
rect 126 37 132 39
rect 95 35 132 37
rect 263 38 308 40
rect 263 36 264 38
rect 266 36 305 38
rect 307 36 308 38
rect 41 30 59 32
rect 41 28 53 30
rect 55 28 59 30
rect 41 26 59 28
rect -62 0 12 5
rect -62 -53 -57 0
rect 47 -11 53 26
rect 80 -2 85 35
rect 263 34 308 36
rect 143 30 171 32
rect 143 28 148 30
rect 150 28 168 30
rect 170 28 171 30
rect 143 26 171 28
rect 215 29 276 30
rect 215 27 216 29
rect 218 27 273 29
rect 275 27 276 29
rect 215 26 276 27
rect 80 -6 220 -2
rect 47 -15 172 -11
rect -52 -20 139 -19
rect -52 -22 -50 -20
rect -48 -22 39 -20
rect 41 -22 132 -20
rect 134 -22 136 -20
rect 138 -22 139 -20
rect -52 -23 139 -22
rect 168 -20 172 -15
rect 216 -17 220 -6
rect 216 -19 217 -17
rect 219 -19 220 -17
rect 216 -20 220 -19
rect 168 -22 169 -20
rect 171 -22 172 -20
rect 168 -24 172 -22
rect 240 -21 292 -20
rect 240 -23 241 -21
rect 243 -23 292 -21
rect 240 -24 292 -23
rect 288 -26 289 -24
rect 291 -26 292 -24
rect 288 -27 292 -26
rect 95 -29 284 -28
rect -31 -31 10 -30
rect -31 -33 -29 -31
rect -27 -33 7 -31
rect 9 -33 10 -31
rect 95 -31 96 -29
rect 98 -31 281 -29
rect 283 -31 284 -29
rect 95 -32 284 -31
rect 303 -29 308 34
rect 303 -31 304 -29
rect 306 -31 308 -29
rect -31 -34 10 -33
rect 303 -36 308 -31
rect 127 -37 161 -36
rect 127 -39 128 -37
rect 130 -39 158 -37
rect 160 -39 161 -37
rect 127 -40 161 -39
rect 260 -37 308 -36
rect 260 -39 261 -37
rect 263 -39 308 -37
rect 260 -40 308 -39
rect -62 -55 -60 -53
rect -58 -55 -57 -53
rect -62 -57 -57 -55
<< alu3 >>
rect 246 46 250 47
rect 246 44 247 46
rect 249 44 250 46
rect 246 5 250 44
rect 131 1 250 5
rect 131 -20 135 1
rect 131 -22 132 -20
rect 134 -22 135 -20
rect 131 -23 135 -22
<< alu4 >>
rect 272 27 276 31
<< ptie >>
rect 9 11 35 13
rect 9 9 11 11
rect 13 9 31 11
rect 33 9 35 11
rect 9 7 35 9
rect 232 12 266 14
rect 232 10 234 12
rect 236 10 262 12
rect 264 10 266 12
rect 232 8 266 10
rect 273 12 279 14
rect 273 10 275 12
rect 277 10 279 12
rect 273 8 279 10
rect 7 -3 13 -1
rect 7 -5 9 -3
rect 11 -5 13 -3
rect 7 -7 13 -5
rect 289 -3 307 -1
rect 289 -5 291 -3
rect 293 -5 303 -3
rect 305 -5 307 -3
rect 289 -7 307 -5
<< ntie >>
rect 40 72 46 74
rect 40 70 42 72
rect 44 70 46 72
rect 40 68 46 70
rect 156 72 162 74
rect 156 70 158 72
rect 160 70 162 72
rect 156 68 162 70
rect 220 72 226 74
rect 220 70 222 72
rect 224 70 226 72
rect 220 68 226 70
rect 232 72 238 74
rect 232 70 234 72
rect 236 70 238 72
rect 273 72 307 74
rect 232 68 238 70
rect 273 70 275 72
rect 277 70 289 72
rect 291 70 303 72
rect 305 70 307 72
rect 273 68 307 70
rect -61 -63 -55 -61
rect -61 -65 -59 -63
rect -57 -65 -55 -63
rect -61 -67 -55 -65
rect 7 -63 13 -61
rect 7 -65 9 -63
rect 11 -65 13 -63
rect 7 -67 13 -65
rect 289 -63 307 -61
rect 289 -65 291 -63
rect 293 -65 303 -63
rect 305 -65 307 -63
rect 289 -67 307 -65
<< nmos >>
rect 16 23 18 29
rect 26 23 28 29
rect 46 17 48 23
rect 56 17 58 23
rect 63 17 65 23
rect 73 17 75 23
rect 80 17 82 23
rect 90 17 92 23
rect 110 17 112 23
rect 120 17 122 23
rect 127 17 129 23
rect 137 17 139 23
rect 144 17 146 23
rect 154 17 156 23
rect 174 17 176 23
rect 184 17 186 23
rect 191 17 193 23
rect 201 17 203 23
rect 208 17 210 23
rect 218 17 220 23
rect 238 20 240 26
rect 248 20 250 26
rect 258 20 260 26
rect 279 20 281 26
rect 291 14 293 23
rect 298 14 300 23
rect -55 -16 -53 -10
rect -45 -16 -43 -10
rect -38 -16 -36 -10
rect -28 -16 -26 -10
rect -21 -16 -19 -10
rect -11 -16 -9 -10
rect 13 -24 15 -15
rect 54 -18 56 -4
rect 23 -24 25 -18
rect 33 -24 35 -18
rect 65 -24 67 -4
rect 72 -24 74 -4
rect 92 -24 94 -10
rect 102 -24 104 -10
rect 112 -17 114 -7
rect 122 -17 124 -4
rect 143 -18 145 -4
rect 154 -24 156 -4
rect 161 -24 163 -4
rect 181 -24 183 -10
rect 191 -24 193 -10
rect 201 -17 203 -7
rect 211 -17 213 -4
rect 231 -18 233 -12
rect 241 -18 243 -10
rect 248 -18 250 -10
rect 258 -18 260 -10
rect 265 -18 267 -10
rect 275 -19 277 -10
rect 295 -24 297 -15
<< pmos >>
rect 18 50 20 70
rect 25 50 27 70
rect 56 51 58 63
rect 63 51 65 63
rect 73 51 75 63
rect 80 51 82 63
rect 90 51 92 63
rect 110 51 112 63
rect 120 51 122 63
rect 127 51 129 63
rect 137 51 139 63
rect 144 51 146 63
rect 46 43 48 49
rect 174 51 176 63
rect 184 51 186 63
rect 191 51 193 63
rect 201 51 203 63
rect 208 51 210 63
rect 154 43 156 49
rect 238 50 240 62
rect 251 53 253 71
rect 258 53 260 71
rect 218 43 220 49
rect 279 43 281 55
rect 289 43 291 53
rect 299 43 301 53
rect -55 -42 -53 -36
rect -45 -56 -43 -44
rect -38 -56 -36 -44
rect -28 -56 -26 -44
rect -21 -56 -19 -44
rect -11 -56 -9 -44
rect 13 -54 15 -36
rect 26 -64 28 -43
rect 33 -64 35 -43
rect 54 -64 56 -36
rect 64 -64 66 -36
rect 74 -64 76 -36
rect 92 -61 94 -36
rect 99 -61 101 -36
rect 109 -52 111 -39
rect 122 -64 124 -39
rect 143 -64 145 -36
rect 153 -64 155 -36
rect 163 -64 165 -36
rect 181 -61 183 -36
rect 188 -61 190 -36
rect 198 -52 200 -39
rect 211 -64 213 -39
rect 231 -44 233 -36
rect 241 -64 243 -48
rect 248 -64 250 -48
rect 258 -64 260 -48
rect 265 -64 267 -48
rect 275 -64 277 -46
rect 295 -54 297 -36
<< polyct0 >>
rect 64 44 66 46
rect 71 28 73 30
rect 136 44 138 46
rect 89 28 91 30
rect 111 28 113 30
rect 129 28 131 30
rect 200 44 202 46
rect 175 28 177 30
rect 193 28 195 30
rect 240 37 242 39
rect 281 36 283 38
rect -30 -23 -28 -21
rect -12 -23 -10 -21
rect -37 -39 -35 -37
rect 15 -31 17 -29
rect 54 -31 56 -29
rect 64 -31 66 -29
rect 120 -24 122 -22
rect 114 -34 116 -32
rect 143 -31 145 -29
rect 153 -31 155 -29
rect 209 -24 211 -22
rect 203 -34 205 -32
rect 256 -25 258 -23
rect 274 -26 276 -24
rect 249 -41 251 -39
<< polyct1 >>
rect 41 54 43 56
rect 17 43 19 45
rect 159 54 161 56
rect 27 34 29 36
rect 54 36 56 38
rect 81 38 83 40
rect 119 38 121 40
rect 223 54 225 56
rect 146 36 148 38
rect 183 38 185 40
rect 291 60 293 62
rect 210 36 212 38
rect 250 44 252 46
rect 260 36 262 38
rect 300 28 302 30
rect -47 -31 -45 -29
rect -20 -33 -18 -31
rect 25 -31 27 -29
rect -60 -49 -58 -47
rect 74 -31 76 -29
rect 81 -31 83 -29
rect 100 -31 102 -29
rect 35 -38 37 -36
rect 163 -31 165 -29
rect 170 -31 172 -29
rect 189 -31 191 -29
rect 239 -31 241 -29
rect 266 -36 268 -34
rect 297 -31 299 -29
rect 226 -51 228 -49
<< ndifct0 >>
rect 10 25 12 27
rect 31 25 33 27
rect 41 19 43 21
rect 51 19 53 21
rect 68 19 70 21
rect 85 19 87 21
rect 115 19 117 21
rect 132 19 134 21
rect 149 19 151 21
rect 159 19 161 21
rect 179 19 181 21
rect 196 19 198 21
rect 213 19 215 21
rect 223 19 225 21
rect 243 22 245 24
rect 253 22 255 24
rect 263 22 265 24
rect 303 19 305 21
rect 19 -9 21 -7
rect -60 -14 -58 -12
rect -50 -14 -48 -12
rect -33 -14 -31 -12
rect -16 -14 -14 -12
rect 38 -9 40 -7
rect 60 -8 62 -6
rect 28 -22 30 -20
rect 77 -15 79 -13
rect 87 -15 89 -13
rect 87 -22 89 -20
rect 97 -22 99 -20
rect 107 -14 109 -12
rect 117 -11 119 -9
rect 149 -8 151 -6
rect 166 -15 168 -13
rect 176 -15 178 -13
rect 176 -22 178 -20
rect 186 -22 188 -20
rect 196 -14 198 -12
rect 206 -11 208 -9
rect 226 -16 228 -14
rect 236 -16 238 -14
rect 253 -14 255 -12
rect 270 -14 272 -12
rect 304 -19 306 -17
<< ndifct1 >>
rect 21 25 23 27
rect 95 19 97 21
rect 105 19 107 21
rect 169 19 171 21
rect 233 22 235 24
rect 274 22 276 24
rect 285 10 287 12
rect -6 -14 -4 -12
rect 8 -22 10 -20
rect 49 -15 51 -13
rect 127 -15 129 -13
rect 138 -15 140 -13
rect 216 -15 218 -13
rect 280 -17 282 -15
rect 290 -22 292 -20
<< ntiect1 >>
rect 42 70 44 72
rect 158 70 160 72
rect 222 70 224 72
rect 234 70 236 72
rect 275 70 277 72
rect 289 70 291 72
rect 303 70 305 72
rect -59 -65 -57 -63
rect 9 -65 11 -63
rect 291 -65 293 -63
rect 303 -65 305 -63
<< ptiect1 >>
rect 11 9 13 11
rect 31 9 33 11
rect 234 10 236 12
rect 262 10 264 12
rect 275 10 277 12
rect 9 -5 11 -3
rect 291 -5 293 -3
rect 303 -5 305 -3
<< pdifct0 >>
rect 32 66 34 68
rect 245 67 247 69
rect 32 59 34 61
rect 51 59 53 61
rect 68 53 70 55
rect 85 59 87 61
rect 115 59 117 61
rect 132 53 134 55
rect 149 59 151 61
rect 41 45 43 47
rect 179 59 181 61
rect 196 53 198 55
rect 213 59 215 61
rect 159 45 161 47
rect 263 60 265 62
rect 223 45 225 47
rect 284 45 286 47
rect 294 45 296 47
rect 304 49 306 51
rect -60 -40 -58 -38
rect -50 -54 -48 -52
rect -33 -48 -31 -46
rect -16 -54 -14 -52
rect 19 -62 21 -60
rect 38 -55 40 -53
rect 59 -55 61 -53
rect 59 -62 61 -60
rect 69 -47 71 -45
rect 69 -54 71 -52
rect 81 -55 83 -53
rect 81 -62 83 -60
rect 104 -43 106 -41
rect 116 -62 118 -60
rect 148 -55 150 -53
rect 148 -62 150 -60
rect 158 -47 160 -45
rect 158 -54 160 -52
rect 170 -55 172 -53
rect 170 -62 172 -60
rect 193 -43 195 -41
rect 205 -62 207 -60
rect 226 -40 228 -38
rect 236 -62 238 -60
rect 253 -52 255 -50
rect 270 -62 272 -60
rect 301 -55 303 -53
<< pdifct1 >>
rect 13 60 15 62
rect 95 53 97 55
rect 105 53 107 55
rect 169 53 171 55
rect 233 58 235 60
rect 274 45 276 47
rect -6 -48 -4 -46
rect 8 -45 10 -43
rect 8 -52 10 -50
rect 49 -40 51 -38
rect 49 -47 51 -45
rect 127 -43 129 -41
rect 127 -50 129 -48
rect 138 -40 140 -38
rect 138 -47 140 -45
rect 216 -43 218 -41
rect 216 -50 218 -48
rect 290 -40 292 -38
rect 290 -47 292 -45
rect 280 -55 282 -53
<< alu0 >>
rect 31 66 32 68
rect 34 66 35 68
rect 31 61 35 66
rect 31 59 32 61
rect 34 59 35 61
rect 31 57 35 59
rect 49 61 55 69
rect 49 59 51 61
rect 53 59 55 61
rect 49 58 55 59
rect 83 61 89 69
rect 83 59 85 61
rect 87 59 89 61
rect 83 58 89 59
rect 113 61 119 69
rect 113 59 115 61
rect 117 59 119 61
rect 113 58 119 59
rect 147 61 153 69
rect 147 59 149 61
rect 151 59 153 61
rect 147 58 153 59
rect 177 61 183 69
rect 177 59 179 61
rect 181 59 183 61
rect 177 58 183 59
rect 211 61 217 69
rect 243 67 245 69
rect 247 67 249 69
rect 243 66 249 67
rect 211 59 213 61
rect 215 59 217 61
rect 211 58 217 59
rect 66 55 72 56
rect 66 53 68 55
rect 70 53 83 55
rect 66 51 83 53
rect 79 48 83 51
rect 39 47 67 48
rect 39 45 41 47
rect 43 46 67 47
rect 43 45 64 46
rect 39 44 64 45
rect 66 44 67 46
rect 9 27 13 29
rect 9 25 10 27
rect 12 25 13 27
rect 9 13 13 25
rect 30 27 35 29
rect 30 25 31 27
rect 33 25 35 27
rect 30 23 35 25
rect 31 13 35 23
rect 39 22 43 44
rect 63 32 67 44
rect 79 44 92 48
rect 63 30 74 32
rect 88 30 92 44
rect 63 28 71 30
rect 73 28 74 30
rect 63 26 74 28
rect 77 28 89 30
rect 91 28 92 30
rect 77 26 92 28
rect 77 22 81 26
rect 39 21 45 22
rect 39 19 41 21
rect 43 19 45 21
rect 39 18 45 19
rect 49 21 55 22
rect 49 19 51 21
rect 53 19 55 21
rect 49 13 55 19
rect 66 21 81 22
rect 66 19 68 21
rect 70 19 81 21
rect 66 18 81 19
rect 84 21 88 23
rect 84 19 85 21
rect 87 19 88 21
rect 84 13 88 19
rect 130 55 136 56
rect 119 53 132 55
rect 134 53 136 55
rect 119 51 136 53
rect 194 55 200 56
rect 183 53 196 55
rect 198 53 200 55
rect 183 51 200 53
rect 247 62 267 63
rect 247 60 263 62
rect 265 60 267 62
rect 247 59 267 60
rect 119 48 123 51
rect 110 44 123 48
rect 135 47 163 48
rect 110 30 114 44
rect 135 46 159 47
rect 135 44 136 46
rect 138 45 159 46
rect 161 45 163 47
rect 138 44 163 45
rect 135 32 139 44
rect 128 30 139 32
rect 110 28 111 30
rect 113 28 125 30
rect 110 26 125 28
rect 128 28 129 30
rect 131 28 139 30
rect 128 26 139 28
rect 114 21 118 23
rect 114 19 115 21
rect 117 19 118 21
rect 114 13 118 19
rect 121 22 125 26
rect 159 22 163 44
rect 121 21 136 22
rect 121 19 132 21
rect 134 19 136 21
rect 121 18 136 19
rect 147 21 153 22
rect 147 19 149 21
rect 151 19 153 21
rect 147 13 153 19
rect 157 21 163 22
rect 157 19 159 21
rect 161 19 163 21
rect 157 18 163 19
rect 183 48 187 51
rect 174 44 187 48
rect 199 47 227 48
rect 174 30 178 44
rect 199 46 223 47
rect 199 44 200 46
rect 202 45 223 46
rect 225 45 227 47
rect 202 44 227 45
rect 199 32 203 44
rect 192 30 203 32
rect 174 28 175 30
rect 177 28 189 30
rect 174 26 189 28
rect 192 28 193 30
rect 195 28 203 30
rect 192 26 203 28
rect 178 21 182 23
rect 178 19 179 21
rect 181 19 182 21
rect 178 13 182 19
rect 185 22 189 26
rect 223 22 227 44
rect 185 21 200 22
rect 185 19 196 21
rect 198 19 200 21
rect 185 18 200 19
rect 211 21 217 22
rect 211 19 213 21
rect 215 19 217 21
rect 211 13 217 19
rect 221 21 227 22
rect 221 19 223 21
rect 225 19 227 21
rect 221 18 227 19
rect 235 56 236 59
rect 247 55 251 59
rect 239 51 251 55
rect 239 39 243 51
rect 239 37 240 39
rect 242 37 243 39
rect 239 32 243 37
rect 239 28 256 32
rect 241 24 247 25
rect 241 22 243 24
rect 245 22 247 24
rect 241 13 247 22
rect 252 24 256 28
rect 276 43 277 49
rect 280 48 284 69
rect 303 51 307 69
rect 303 49 304 51
rect 306 49 307 51
rect 280 47 288 48
rect 280 45 284 47
rect 286 45 288 47
rect 280 44 288 45
rect 292 47 298 48
rect 303 47 307 49
rect 292 45 294 47
rect 296 45 298 47
rect 292 39 298 45
rect 279 38 298 39
rect 279 36 281 38
rect 283 36 298 38
rect 279 35 298 36
rect 252 22 253 24
rect 255 22 256 24
rect 252 20 256 22
rect 261 24 267 25
rect 261 22 263 24
rect 265 22 267 24
rect 261 13 267 22
rect 276 24 277 26
rect 288 22 292 35
rect 288 21 307 22
rect 288 19 303 21
rect 305 19 307 21
rect 288 18 307 19
rect -62 -12 -56 -11
rect -62 -14 -60 -12
rect -58 -14 -56 -12
rect -62 -15 -56 -14
rect -52 -12 -46 -6
rect -52 -14 -50 -12
rect -48 -14 -46 -12
rect -52 -15 -46 -14
rect -35 -12 -20 -11
rect -35 -14 -33 -12
rect -31 -14 -20 -12
rect -35 -15 -20 -14
rect -62 -37 -58 -15
rect -24 -19 -20 -15
rect -17 -12 -13 -6
rect 17 -7 23 -6
rect 17 -9 19 -7
rect 21 -9 23 -7
rect 17 -10 23 -9
rect 36 -7 42 -6
rect 36 -9 38 -7
rect 40 -9 42 -7
rect 58 -8 60 -6
rect 62 -8 64 -6
rect 58 -9 64 -8
rect 116 -9 120 -6
rect 147 -8 149 -6
rect 151 -8 153 -6
rect 147 -9 153 -8
rect 205 -9 209 -6
rect 36 -10 42 -9
rect 116 -11 117 -9
rect 119 -11 120 -9
rect 205 -11 206 -9
rect 208 -11 209 -9
rect -17 -14 -16 -12
rect -14 -14 -13 -12
rect -17 -16 -13 -14
rect 86 -12 111 -11
rect -38 -21 -27 -19
rect -38 -23 -30 -21
rect -28 -23 -27 -21
rect -24 -21 -9 -19
rect -24 -23 -12 -21
rect -10 -23 -9 -21
rect -38 -25 -27 -23
rect -38 -37 -34 -25
rect -62 -38 -37 -37
rect -62 -40 -60 -38
rect -58 -39 -37 -38
rect -35 -39 -34 -37
rect -58 -40 -34 -39
rect -13 -37 -9 -23
rect -62 -41 -34 -40
rect -22 -41 -9 -37
rect -22 -44 -18 -41
rect 71 -13 81 -12
rect 71 -15 77 -13
rect 79 -15 81 -13
rect 71 -16 81 -15
rect 86 -13 107 -12
rect 86 -15 87 -13
rect 89 -14 107 -13
rect 109 -14 111 -12
rect 116 -13 120 -11
rect 175 -12 200 -11
rect 89 -15 111 -14
rect -35 -46 -18 -44
rect -35 -48 -33 -46
rect -31 -48 -18 -46
rect -35 -49 -29 -48
rect 14 -20 32 -19
rect 14 -22 28 -20
rect 30 -22 32 -20
rect 14 -23 32 -22
rect 14 -29 18 -23
rect 14 -31 15 -29
rect 17 -31 18 -29
rect -52 -52 -46 -51
rect -52 -54 -50 -52
rect -48 -54 -46 -52
rect -52 -62 -46 -54
rect -18 -52 -12 -51
rect -18 -54 -16 -52
rect -14 -54 -12 -52
rect -18 -62 -12 -54
rect 10 -52 11 -41
rect 14 -44 18 -31
rect 33 -36 39 -35
rect 71 -20 75 -16
rect 55 -24 75 -20
rect 55 -27 59 -24
rect 53 -29 59 -27
rect 53 -31 54 -29
rect 56 -31 59 -29
rect 53 -33 59 -31
rect 14 -48 29 -44
rect 25 -52 29 -48
rect 55 -44 59 -33
rect 63 -29 67 -27
rect 86 -20 90 -15
rect 86 -22 87 -20
rect 89 -22 90 -20
rect 86 -24 90 -22
rect 95 -20 110 -19
rect 95 -22 97 -20
rect 99 -21 110 -20
rect 99 -22 124 -21
rect 95 -23 120 -22
rect 106 -24 120 -23
rect 122 -24 124 -22
rect 106 -25 124 -24
rect 63 -31 64 -29
rect 66 -31 67 -29
rect 63 -36 67 -31
rect 106 -36 110 -25
rect 103 -40 110 -36
rect 113 -32 117 -30
rect 113 -34 114 -32
rect 116 -34 117 -32
rect 103 -41 107 -40
rect 103 -43 104 -41
rect 106 -43 107 -41
rect 55 -45 95 -44
rect 103 -45 107 -43
rect 113 -44 117 -34
rect 55 -47 69 -45
rect 71 -47 95 -45
rect 55 -48 95 -47
rect 111 -48 117 -44
rect 68 -52 72 -48
rect 91 -52 115 -48
rect 160 -13 170 -12
rect 160 -15 166 -13
rect 168 -15 170 -13
rect 160 -16 170 -15
rect 175 -13 196 -12
rect 175 -15 176 -13
rect 178 -14 196 -13
rect 198 -14 200 -12
rect 205 -13 209 -11
rect 178 -15 200 -14
rect 160 -20 164 -16
rect 144 -24 164 -20
rect 144 -27 148 -24
rect 142 -29 148 -27
rect 142 -31 143 -29
rect 145 -31 148 -29
rect 142 -33 148 -31
rect 144 -44 148 -33
rect 152 -29 156 -27
rect 175 -20 179 -15
rect 175 -22 176 -20
rect 178 -22 179 -20
rect 175 -24 179 -22
rect 184 -20 199 -19
rect 184 -22 186 -20
rect 188 -21 199 -20
rect 188 -22 213 -21
rect 184 -23 209 -22
rect 195 -24 209 -23
rect 211 -24 213 -22
rect 195 -25 213 -24
rect 152 -31 153 -29
rect 155 -31 156 -29
rect 152 -36 156 -31
rect 195 -36 199 -25
rect 192 -40 199 -36
rect 202 -32 206 -30
rect 202 -34 203 -32
rect 205 -34 206 -32
rect 192 -41 196 -40
rect 192 -43 193 -41
rect 195 -43 196 -41
rect 144 -45 184 -44
rect 192 -45 196 -43
rect 202 -44 206 -34
rect 144 -47 158 -45
rect 160 -47 184 -45
rect 144 -48 184 -47
rect 200 -48 206 -44
rect 224 -14 230 -13
rect 224 -16 226 -14
rect 228 -16 230 -14
rect 224 -17 230 -16
rect 234 -14 240 -6
rect 234 -16 236 -14
rect 238 -16 240 -14
rect 251 -12 266 -11
rect 251 -14 253 -12
rect 255 -14 266 -12
rect 251 -15 266 -14
rect 234 -17 240 -16
rect 224 -37 228 -17
rect 262 -20 266 -15
rect 269 -12 273 -6
rect 269 -14 270 -12
rect 272 -14 273 -12
rect 269 -16 273 -14
rect 248 -23 259 -21
rect 248 -25 256 -23
rect 258 -25 259 -23
rect 262 -22 276 -20
rect 262 -24 277 -22
rect 248 -27 259 -25
rect 272 -26 274 -24
rect 276 -26 277 -24
rect 248 -37 252 -27
rect 272 -28 277 -26
rect 224 -38 252 -37
rect 224 -40 226 -38
rect 228 -39 252 -38
rect 228 -40 249 -39
rect 224 -41 249 -40
rect 251 -41 252 -39
rect 268 -38 269 -32
rect 248 -43 252 -41
rect 157 -52 161 -48
rect 180 -52 204 -48
rect 25 -53 42 -52
rect 25 -55 38 -53
rect 40 -55 42 -53
rect 25 -56 42 -55
rect 57 -53 63 -52
rect 57 -55 59 -53
rect 61 -55 63 -53
rect 17 -60 23 -59
rect 17 -62 19 -60
rect 21 -62 23 -60
rect 57 -60 63 -55
rect 68 -54 69 -52
rect 71 -54 72 -52
rect 68 -56 72 -54
rect 79 -53 85 -52
rect 79 -55 81 -53
rect 83 -55 85 -53
rect 57 -62 59 -60
rect 61 -62 63 -60
rect 79 -60 85 -55
rect 146 -53 152 -52
rect 146 -55 148 -53
rect 150 -55 152 -53
rect 79 -62 81 -60
rect 83 -62 85 -60
rect 114 -60 120 -59
rect 114 -62 116 -60
rect 118 -62 120 -60
rect 146 -60 152 -55
rect 157 -54 158 -52
rect 160 -54 161 -52
rect 157 -56 161 -54
rect 168 -53 174 -52
rect 168 -55 170 -53
rect 172 -55 174 -53
rect 146 -62 148 -60
rect 150 -62 152 -60
rect 168 -60 174 -55
rect 272 -45 276 -28
rect 260 -49 276 -45
rect 251 -50 264 -49
rect 251 -52 253 -50
rect 255 -52 264 -50
rect 303 -17 307 -6
rect 292 -24 293 -18
rect 303 -19 304 -17
rect 306 -19 307 -17
rect 303 -21 307 -19
rect 292 -43 293 -36
rect 251 -53 264 -52
rect 299 -53 305 -52
rect 299 -55 301 -53
rect 303 -55 305 -53
rect 168 -62 170 -60
rect 172 -62 174 -60
rect 203 -60 209 -59
rect 203 -62 205 -60
rect 207 -62 209 -60
rect 235 -60 239 -58
rect 235 -62 236 -60
rect 238 -62 239 -60
rect 268 -60 274 -59
rect 268 -62 270 -60
rect 272 -62 274 -60
rect 299 -62 305 -55
<< via1 >>
rect 40 59 42 61
rect 160 58 162 60
rect 224 59 226 61
rect 25 52 27 54
rect 9 40 11 42
rect 33 44 35 46
rect 53 28 55 30
rect 76 37 78 39
rect 96 37 98 39
rect 124 37 126 39
rect 148 28 150 30
rect 168 28 170 30
rect 193 40 195 42
rect 216 27 218 29
rect 232 40 234 42
rect 256 53 258 55
rect 264 36 266 38
rect 289 53 291 55
rect 305 36 307 38
rect 273 27 275 29
rect -50 -22 -48 -20
rect -29 -33 -27 -31
rect 39 -22 41 -20
rect 7 -33 9 -31
rect -60 -55 -58 -53
rect 96 -31 98 -29
rect 128 -39 130 -37
rect 136 -22 138 -20
rect 169 -22 171 -20
rect 217 -19 219 -17
rect 158 -39 160 -37
rect 241 -23 243 -21
rect 261 -39 263 -37
rect 281 -31 283 -29
rect 289 -26 291 -24
rect 304 -31 306 -29
<< via2 >>
rect 247 44 249 46
rect 132 -22 134 -20
<< labels >>
rlabel alu1 134 -2 134 -2 5 Vss
rlabel alu1 226 -56 226 -56 5 Binv
rlabel alu1 218 -33 218 -33 5 Sum
rlabel via1 262 -38 262 -38 5 B
rlabel alu1 81 -20 81 -20 5 A
rlabel alu1 134 -66 134 -66 5 Vdd
rlabel alu1 170 -22 170 -22 5 Cin
rlabel alu1 -4 -34 -4 -34 1 COUT
rlabel alu1 -32 -66 -32 -66 2 vdd
rlabel alu1 -32 -2 -32 -2 2 vss
rlabel alu1 69 9 69 9 4 vss
rlabel alu1 69 73 69 73 4 vdd
rlabel alu1 133 9 133 9 6 vss
rlabel alu1 133 73 133 73 6 vdd
rlabel alu1 197 73 197 73 6 vdd
rlabel alu1 197 9 197 9 6 vss
rlabel alu1 290 73 290 73 6 vdd
rlabel alu1 249 9 249 9 6 vss
rlabel alu1 249 73 249 73 6 vdd
rlabel space 229 8 269 76 1 or
rlabel space 271 8 311 76 1 and
rlabel space 32 8 229 76 1 4x1_mux
rlabel alu1 290 9 290 9 6 vss
rlabel space 1 -70 312 6 1 fafs
rlabel space -64 -70 0 6 1 shift_mux
rlabel alu1 22 8 22 8 6 vss
rlabel alu1 22 72 22 72 6 vdd
rlabel ab 7 7 36 76 1 decoder
rlabel alu1 160 63 160 63 1 s1
rlabel alu2 99 60 99 60 1 s0
<< end >>
