magic
tech scmos
timestamp 1760355489
<< ab >>
rect -155 75 -46 147
rect -44 75 -2 147
rect 0 75 63 147
rect 70 77 100 147
rect 101 146 178 147
rect 185 146 291 147
rect 297 146 374 147
rect 101 78 333 146
rect 334 78 374 146
rect 65 75 97 77
rect -33 71 -1 73
rect -310 2 -270 70
rect -269 2 -37 70
rect -310 1 -233 2
rect -227 1 -121 2
rect -114 1 -37 2
rect -36 1 -6 71
rect 1 1 64 73
rect 66 1 108 73
rect 110 1 219 73
<< nwell >>
rect -312 108 376 147
rect -312 107 70 108
rect -4 40 24 41
rect 63 40 376 41
rect -312 1 376 40
<< pwell >>
rect 70 107 376 108
rect -312 67 376 107
rect -312 41 4 67
rect 24 41 376 67
rect -312 40 -4 41
rect 24 40 63 41
<< poly >>
rect -277 141 -275 145
rect -267 141 -265 145
rect -260 141 -258 145
rect -250 141 -248 145
rect -243 141 -241 145
rect -213 141 -211 145
rect -297 131 -295 136
rect -230 128 -224 130
rect -230 126 -228 128
rect -226 126 -224 128
rect -297 110 -295 113
rect -301 108 -295 110
rect -301 106 -299 108
rect -297 106 -295 108
rect -301 104 -295 106
rect -277 105 -275 123
rect -267 115 -265 125
rect -270 113 -264 115
rect -270 111 -268 113
rect -266 111 -264 113
rect -270 109 -264 111
rect -260 110 -258 125
rect -250 120 -248 125
rect -253 118 -247 120
rect -253 116 -251 118
rect -249 116 -247 118
rect -253 114 -247 116
rect -243 110 -241 125
rect -233 124 -224 126
rect -233 121 -231 124
rect -190 138 -188 143
rect -183 138 -181 143
rect -165 141 -163 145
rect -155 141 -153 145
rect -145 141 -143 145
rect -124 141 -122 145
rect -200 129 -198 134
rect -297 101 -295 104
rect -278 103 -272 105
rect -278 101 -276 103
rect -274 101 -272 103
rect -278 99 -272 101
rect -277 96 -275 99
rect -297 87 -295 92
rect -267 95 -265 109
rect -260 108 -248 110
rect -260 102 -254 104
rect -260 100 -258 102
rect -256 100 -254 102
rect -260 98 -254 100
rect -260 95 -258 98
rect -250 95 -248 108
rect -243 108 -237 110
rect -243 106 -241 108
rect -239 106 -237 108
rect -243 104 -237 106
rect -243 95 -241 104
rect -233 95 -231 113
rect -213 103 -211 116
rect -200 113 -198 116
rect -101 138 -99 143
rect -94 138 -92 143
rect -76 141 -74 145
rect -66 141 -64 145
rect -56 141 -54 145
rect -35 141 -33 145
rect -28 141 -26 145
rect -111 129 -109 134
rect -207 111 -198 113
rect -207 109 -205 111
rect -203 109 -201 111
rect -190 110 -188 113
rect -183 110 -181 113
rect -165 110 -163 113
rect -155 110 -153 113
rect -145 110 -143 113
rect -207 107 -201 109
rect -213 101 -207 103
rect -213 99 -211 101
rect -209 99 -207 101
rect -213 97 -207 99
rect -213 94 -211 97
rect -203 94 -201 107
rect -193 108 -187 110
rect -193 106 -191 108
rect -189 106 -187 108
rect -193 104 -187 106
rect -183 108 -161 110
rect -183 106 -172 108
rect -170 106 -165 108
rect -163 106 -161 108
rect -183 104 -161 106
rect -157 108 -151 110
rect -157 106 -155 108
rect -153 106 -151 108
rect -157 104 -151 106
rect -147 108 -141 110
rect -147 106 -145 108
rect -143 106 -141 108
rect -147 104 -141 106
rect -193 101 -191 104
rect -183 101 -181 104
rect -163 101 -161 104
rect -156 101 -154 104
rect -277 82 -275 87
rect -267 82 -265 87
rect -260 82 -258 87
rect -250 79 -248 87
rect -243 83 -241 87
rect -233 79 -231 89
rect -250 77 -231 79
rect -213 77 -211 81
rect -203 79 -201 84
rect -193 82 -191 87
rect -183 82 -181 87
rect -145 95 -143 104
rect -124 103 -122 116
rect -111 113 -109 116
rect 82 141 84 145
rect 89 141 91 145
rect -15 131 -13 136
rect 9 133 11 138
rect 19 133 21 138
rect 26 133 28 138
rect 36 133 38 138
rect 43 133 45 138
rect -35 117 -33 120
rect -39 115 -33 117
rect -39 113 -37 115
rect -35 113 -33 115
rect -118 111 -109 113
rect -118 109 -116 111
rect -114 109 -112 111
rect -101 110 -99 113
rect -94 110 -92 113
rect -76 110 -74 113
rect -66 110 -64 113
rect -56 110 -54 113
rect -39 111 -33 113
rect -118 107 -112 109
rect -124 101 -118 103
rect -124 99 -122 101
rect -120 99 -118 101
rect -124 97 -118 99
rect -124 94 -122 97
rect -114 94 -112 107
rect -104 108 -98 110
rect -104 106 -102 108
rect -100 106 -98 108
rect -104 104 -98 106
rect -94 108 -72 110
rect -94 106 -83 108
rect -81 106 -76 108
rect -74 106 -72 108
rect -94 104 -72 106
rect -68 108 -62 110
rect -68 106 -66 108
rect -64 106 -62 108
rect -68 104 -62 106
rect -58 108 -52 110
rect -58 106 -56 108
rect -54 106 -52 108
rect -58 104 -52 106
rect -104 101 -102 104
rect -94 101 -92 104
rect -74 101 -72 104
rect -67 101 -65 104
rect -163 77 -161 81
rect -156 77 -154 81
rect -145 77 -143 81
rect -124 77 -122 81
rect -114 79 -112 84
rect -104 82 -102 87
rect -94 82 -92 87
rect -56 95 -54 104
rect -35 101 -33 111
rect -28 110 -26 120
rect 56 126 62 128
rect 56 124 58 126
rect 60 124 62 126
rect -15 110 -13 113
rect -29 108 -23 110
rect -29 106 -27 108
rect -25 106 -23 108
rect -29 104 -23 106
rect -19 108 -13 110
rect -19 106 -17 108
rect -15 106 -13 108
rect -19 104 -13 106
rect -25 101 -23 104
rect -15 101 -13 104
rect 9 102 11 121
rect 19 112 21 121
rect 16 110 22 112
rect 16 108 18 110
rect 20 108 22 110
rect 16 106 22 108
rect 26 108 28 121
rect 36 118 38 121
rect 33 116 39 118
rect 33 114 35 116
rect 37 114 39 116
rect 33 112 39 114
rect 43 110 45 121
rect 53 122 62 124
rect 53 119 55 122
rect 315 142 317 146
rect 322 142 324 146
rect 120 134 122 139
rect 127 134 129 139
rect 137 134 139 139
rect 144 134 146 139
rect 154 134 156 139
rect 174 134 176 139
rect 184 134 186 139
rect 191 134 193 139
rect 201 134 203 139
rect 208 134 210 139
rect 238 134 240 139
rect 248 134 250 139
rect 255 134 257 139
rect 265 134 267 139
rect 272 134 274 139
rect 103 127 109 129
rect 103 125 105 127
rect 107 125 109 127
rect 103 123 112 125
rect 82 118 84 121
rect 79 116 85 118
rect 79 114 81 116
rect 83 114 85 116
rect 43 108 49 110
rect 26 106 38 108
rect -35 90 -33 95
rect -25 90 -23 95
rect 8 100 14 102
rect 8 98 10 100
rect 12 98 14 100
rect 8 96 14 98
rect 9 93 11 96
rect 19 93 21 106
rect 26 100 32 102
rect 26 98 28 100
rect 30 98 32 100
rect 26 96 32 98
rect 26 93 28 96
rect 36 93 38 106
rect 43 106 45 108
rect 47 106 49 108
rect 43 104 49 106
rect 43 93 45 104
rect 53 93 55 113
rect 79 112 85 114
rect 80 100 82 112
rect 89 109 91 121
rect 110 120 112 123
rect 221 127 227 129
rect 221 125 223 127
rect 225 125 227 127
rect 89 107 95 109
rect 89 105 91 107
rect 93 105 95 107
rect 89 103 95 105
rect 90 100 92 103
rect 110 94 112 114
rect 120 111 122 122
rect 127 119 129 122
rect 126 117 132 119
rect 126 115 128 117
rect 130 115 132 117
rect 126 113 132 115
rect 116 109 122 111
rect 137 109 139 122
rect 144 113 146 122
rect 116 107 118 109
rect 120 107 122 109
rect 116 105 122 107
rect 120 94 122 105
rect 127 107 139 109
rect 143 111 149 113
rect 143 109 145 111
rect 147 109 149 111
rect 143 107 149 109
rect 127 94 129 107
rect 133 101 139 103
rect 133 99 135 101
rect 137 99 139 101
rect 133 97 139 99
rect 137 94 139 97
rect 144 94 146 107
rect 154 103 156 122
rect 174 103 176 122
rect 184 113 186 122
rect 181 111 187 113
rect 181 109 183 111
rect 185 109 187 111
rect 181 107 187 109
rect 191 109 193 122
rect 201 119 203 122
rect 198 117 204 119
rect 198 115 200 117
rect 202 115 204 117
rect 198 113 204 115
rect 208 111 210 122
rect 218 123 227 125
rect 218 120 220 123
rect 302 133 304 137
rect 285 127 291 129
rect 285 125 287 127
rect 289 125 291 127
rect 208 109 214 111
rect 191 107 203 109
rect 151 101 157 103
rect 151 99 153 101
rect 155 99 157 101
rect 151 97 157 99
rect 173 101 179 103
rect 173 99 175 101
rect 177 99 179 101
rect 173 97 179 99
rect 154 94 156 97
rect 174 94 176 97
rect 184 94 186 107
rect 191 101 197 103
rect 191 99 193 101
rect 195 99 197 101
rect 191 97 197 99
rect 191 94 193 97
rect 201 94 203 107
rect 208 107 210 109
rect 212 107 214 109
rect 208 105 214 107
rect 208 94 210 105
rect 218 94 220 114
rect 238 103 240 122
rect 248 113 250 122
rect 245 111 251 113
rect 245 109 247 111
rect 249 109 251 111
rect 245 107 251 109
rect 255 109 257 122
rect 265 119 267 122
rect 262 117 268 119
rect 262 115 264 117
rect 266 115 268 117
rect 262 113 268 115
rect 272 111 274 122
rect 282 123 291 125
rect 282 120 284 123
rect 353 133 359 135
rect 353 131 355 133
rect 357 131 359 133
rect 343 126 345 131
rect 353 129 359 131
rect 272 109 278 111
rect 255 107 267 109
rect 237 101 243 103
rect 237 99 239 101
rect 241 99 243 101
rect 237 97 243 99
rect 238 94 240 97
rect 248 94 250 107
rect 255 101 261 103
rect 255 99 257 101
rect 259 99 261 101
rect 255 97 261 99
rect 255 94 257 97
rect 265 94 267 107
rect 272 107 274 109
rect 276 107 278 109
rect 272 105 278 107
rect 272 94 274 105
rect 282 94 284 114
rect 302 112 304 121
rect 315 119 317 124
rect 312 117 318 119
rect 312 115 314 117
rect 316 115 318 117
rect 312 113 318 115
rect 302 110 308 112
rect 302 108 304 110
rect 306 108 308 110
rect 302 106 308 108
rect 302 97 304 106
rect 312 97 314 113
rect 322 111 324 124
rect 353 124 355 129
rect 363 124 365 129
rect 343 111 345 114
rect 353 111 355 114
rect 322 109 328 111
rect 322 107 324 109
rect 326 107 328 109
rect 322 105 328 107
rect 343 109 349 111
rect 343 107 345 109
rect 347 107 349 109
rect 353 108 357 111
rect 343 105 349 107
rect 322 97 324 105
rect 343 97 345 105
rect -15 87 -13 92
rect 80 89 82 94
rect 90 89 92 94
rect 355 94 357 108
rect 363 103 365 114
rect 362 101 368 103
rect 362 99 364 101
rect 366 99 368 101
rect 362 97 368 99
rect 362 94 364 97
rect 9 82 11 87
rect 19 82 21 87
rect 26 82 28 87
rect -74 77 -72 81
rect -67 77 -65 81
rect -56 77 -54 81
rect 36 79 38 87
rect 43 83 45 87
rect 53 79 55 87
rect 36 77 55 79
rect 110 80 112 88
rect 120 84 122 88
rect 127 80 129 88
rect 137 83 139 88
rect 144 83 146 88
rect 154 83 156 88
rect 174 83 176 88
rect 184 83 186 88
rect 191 83 193 88
rect 110 78 129 80
rect 201 80 203 88
rect 208 84 210 88
rect 218 80 220 88
rect 238 83 240 88
rect 248 83 250 88
rect 255 83 257 88
rect 201 78 220 80
rect 265 80 267 88
rect 272 84 274 88
rect 282 80 284 88
rect 302 87 304 91
rect 312 87 314 91
rect 322 87 324 91
rect 343 87 345 91
rect 265 78 284 80
rect 355 80 357 85
rect 362 80 364 85
rect -300 63 -298 68
rect -293 63 -291 68
rect -220 68 -201 70
rect -281 57 -279 61
rect -260 57 -258 61
rect -250 57 -248 61
rect -240 57 -238 61
rect -220 60 -218 68
rect -210 60 -208 64
rect -203 60 -201 68
rect -156 68 -137 70
rect -193 60 -191 65
rect -186 60 -184 65
rect -176 60 -174 65
rect -156 60 -154 68
rect -146 60 -144 64
rect -139 60 -137 68
rect -65 68 -46 70
rect -129 60 -127 65
rect -122 60 -120 65
rect -112 60 -110 65
rect -92 60 -90 65
rect -82 60 -80 65
rect -75 60 -73 65
rect -65 60 -63 68
rect -58 60 -56 64
rect -48 60 -46 68
rect 9 69 28 71
rect 9 61 11 69
rect 19 61 21 65
rect 26 61 28 69
rect 118 67 120 71
rect 129 67 131 71
rect 136 67 138 71
rect 36 61 38 66
rect 43 61 45 66
rect 53 61 55 66
rect -300 51 -298 54
rect -304 49 -298 51
rect -304 47 -302 49
rect -300 47 -298 49
rect -304 45 -298 47
rect -301 34 -299 45
rect -293 40 -291 54
rect -28 54 -26 59
rect -18 54 -16 59
rect 77 56 79 61
rect -281 43 -279 51
rect -260 43 -258 51
rect -285 41 -279 43
rect -293 37 -289 40
rect -285 39 -283 41
rect -281 39 -279 41
rect -285 37 -279 39
rect -264 41 -258 43
rect -264 39 -262 41
rect -260 39 -258 41
rect -264 37 -258 39
rect -291 34 -289 37
rect -281 34 -279 37
rect -301 19 -299 24
rect -291 19 -289 24
rect -260 24 -258 37
rect -250 35 -248 51
rect -240 42 -238 51
rect -244 40 -238 42
rect -244 38 -242 40
rect -240 38 -238 40
rect -244 36 -238 38
rect -254 33 -248 35
rect -254 31 -252 33
rect -250 31 -248 33
rect -254 29 -248 31
rect -253 24 -251 29
rect -240 27 -238 36
rect -220 34 -218 54
rect -210 43 -208 54
rect -214 41 -208 43
rect -214 39 -212 41
rect -210 39 -208 41
rect -203 41 -201 54
rect -193 51 -191 54
rect -197 49 -191 51
rect -197 47 -195 49
rect -193 47 -191 49
rect -197 45 -191 47
rect -186 41 -184 54
rect -176 51 -174 54
rect -179 49 -173 51
rect -179 47 -177 49
rect -175 47 -173 49
rect -179 45 -173 47
rect -203 39 -191 41
rect -214 37 -208 39
rect -295 17 -289 19
rect -281 17 -279 22
rect -295 15 -293 17
rect -291 15 -289 17
rect -295 13 -289 15
rect -220 25 -218 28
rect -227 23 -218 25
rect -210 26 -208 37
rect -204 33 -198 35
rect -204 31 -202 33
rect -200 31 -198 33
rect -204 29 -198 31
rect -203 26 -201 29
rect -193 26 -191 39
rect -187 39 -181 41
rect -187 37 -185 39
rect -183 37 -181 39
rect -187 35 -181 37
rect -186 26 -184 35
rect -176 26 -174 45
rect -156 34 -154 54
rect -146 43 -144 54
rect -150 41 -144 43
rect -150 39 -148 41
rect -146 39 -144 41
rect -139 41 -137 54
rect -129 51 -127 54
rect -133 49 -127 51
rect -133 47 -131 49
rect -129 47 -127 49
rect -133 45 -127 47
rect -122 41 -120 54
rect -112 51 -110 54
rect -92 51 -90 54
rect -115 49 -109 51
rect -115 47 -113 49
rect -111 47 -109 49
rect -115 45 -109 47
rect -93 49 -87 51
rect -93 47 -91 49
rect -89 47 -87 49
rect -93 45 -87 47
rect -139 39 -127 41
rect -150 37 -144 39
rect -227 21 -225 23
rect -223 21 -221 23
rect -227 19 -221 21
rect -240 11 -238 15
rect -156 25 -154 28
rect -163 23 -154 25
rect -146 26 -144 37
rect -140 33 -134 35
rect -140 31 -138 33
rect -136 31 -134 33
rect -140 29 -134 31
rect -139 26 -137 29
rect -129 26 -127 39
rect -123 39 -117 41
rect -123 37 -121 39
rect -119 37 -117 39
rect -123 35 -117 37
rect -122 26 -120 35
rect -112 26 -110 45
rect -92 26 -90 45
rect -82 41 -80 54
rect -75 51 -73 54
rect -75 49 -69 51
rect -75 47 -73 49
rect -71 47 -69 49
rect -75 45 -69 47
rect -65 41 -63 54
rect -85 39 -79 41
rect -85 37 -83 39
rect -81 37 -79 39
rect -85 35 -79 37
rect -75 39 -63 41
rect -58 43 -56 54
rect -58 41 -52 43
rect -58 39 -56 41
rect -54 39 -52 41
rect -82 26 -80 35
rect -75 26 -73 39
rect -58 37 -52 39
rect -68 33 -62 35
rect -68 31 -66 33
rect -64 31 -62 33
rect -68 29 -62 31
rect -65 26 -63 29
rect -58 26 -56 37
rect -48 34 -46 54
rect -28 45 -26 48
rect -31 43 -25 45
rect -31 41 -29 43
rect -27 41 -25 43
rect -31 39 -25 41
rect -163 21 -161 23
rect -159 21 -157 23
rect -163 19 -157 21
rect -48 25 -46 28
rect -27 27 -25 39
rect -18 36 -16 48
rect -21 34 -15 36
rect 9 35 11 55
rect 19 44 21 55
rect 15 42 21 44
rect 15 40 17 42
rect 19 40 21 42
rect 26 42 28 55
rect 36 52 38 55
rect 32 50 38 52
rect 32 48 34 50
rect 36 48 38 50
rect 32 46 38 48
rect 43 42 45 55
rect 53 52 55 55
rect 50 50 56 52
rect 50 48 52 50
rect 54 48 56 50
rect 50 46 56 48
rect 87 53 89 58
rect 97 53 99 58
rect 26 40 38 42
rect 15 38 21 40
rect -21 32 -19 34
rect -17 32 -15 34
rect -21 30 -15 32
rect -20 27 -18 30
rect -48 23 -39 25
rect -45 21 -43 23
rect -41 21 -39 23
rect -45 19 -39 21
rect -210 9 -208 14
rect -203 9 -201 14
rect -193 9 -191 14
rect -186 9 -184 14
rect -176 9 -174 14
rect -146 9 -144 14
rect -139 9 -137 14
rect -129 9 -127 14
rect -122 9 -120 14
rect -112 9 -110 14
rect -92 9 -90 14
rect -82 9 -80 14
rect -75 9 -73 14
rect -65 9 -63 14
rect -58 9 -56 14
rect -260 2 -258 6
rect -253 2 -251 6
rect 9 26 11 29
rect 2 24 11 26
rect 19 27 21 38
rect 25 34 31 36
rect 25 32 27 34
rect 29 32 31 34
rect 25 30 31 32
rect 26 27 28 30
rect 36 27 38 40
rect 42 40 48 42
rect 42 38 44 40
rect 46 38 48 40
rect 42 36 48 38
rect 43 27 45 36
rect 53 27 55 46
rect 77 44 79 47
rect 87 44 89 47
rect 77 42 83 44
rect 77 40 79 42
rect 81 40 83 42
rect 77 38 83 40
rect 87 42 93 44
rect 87 40 89 42
rect 91 40 93 42
rect 87 38 93 40
rect 77 35 79 38
rect 2 22 4 24
rect 6 22 8 24
rect 2 20 8 22
rect 90 28 92 38
rect 97 37 99 47
rect 118 44 120 53
rect 156 61 158 66
rect 166 61 168 66
rect 176 64 178 69
rect 186 67 188 71
rect 207 67 209 71
rect 218 67 220 71
rect 225 67 227 71
rect 129 44 131 47
rect 136 44 138 47
rect 156 44 158 47
rect 166 44 168 47
rect 116 42 122 44
rect 116 40 118 42
rect 120 40 122 42
rect 116 38 122 40
rect 126 42 132 44
rect 126 40 128 42
rect 130 40 132 42
rect 126 38 132 40
rect 136 42 158 44
rect 136 40 138 42
rect 140 40 145 42
rect 147 40 158 42
rect 136 38 158 40
rect 162 42 168 44
rect 162 40 164 42
rect 166 40 168 42
rect 162 38 168 40
rect 176 41 178 54
rect 186 51 188 54
rect 182 49 188 51
rect 182 47 184 49
rect 186 47 188 49
rect 182 45 188 47
rect 176 39 182 41
rect 97 35 103 37
rect 118 35 120 38
rect 128 35 130 38
rect 138 35 140 38
rect 156 35 158 38
rect 163 35 165 38
rect 176 37 178 39
rect 180 37 182 39
rect 173 35 182 37
rect 97 33 99 35
rect 101 33 103 35
rect 97 31 103 33
rect 97 28 99 31
rect 19 10 21 15
rect 26 10 28 15
rect 36 10 38 15
rect 43 10 45 15
rect 53 10 55 15
rect 77 12 79 17
rect -27 3 -25 7
rect -20 3 -18 7
rect 173 32 175 35
rect 186 32 188 45
rect 207 44 209 53
rect 245 61 247 66
rect 255 61 257 66
rect 265 64 267 69
rect 275 67 277 71
rect 295 69 314 71
rect 295 59 297 69
rect 305 61 307 65
rect 312 61 314 69
rect 322 61 324 66
rect 329 61 331 66
rect 339 61 341 66
rect 218 44 220 47
rect 225 44 227 47
rect 245 44 247 47
rect 255 44 257 47
rect 205 42 211 44
rect 205 40 207 42
rect 209 40 211 42
rect 205 38 211 40
rect 215 42 221 44
rect 215 40 217 42
rect 219 40 221 42
rect 215 38 221 40
rect 225 42 247 44
rect 225 40 227 42
rect 229 40 234 42
rect 236 40 247 42
rect 225 38 247 40
rect 251 42 257 44
rect 251 40 253 42
rect 255 40 257 42
rect 251 38 257 40
rect 265 41 267 54
rect 275 51 277 54
rect 271 49 277 51
rect 271 47 273 49
rect 275 47 277 49
rect 271 45 277 47
rect 265 39 271 41
rect 207 35 209 38
rect 217 35 219 38
rect 227 35 229 38
rect 245 35 247 38
rect 252 35 254 38
rect 265 37 267 39
rect 269 37 271 39
rect 262 35 271 37
rect 173 14 175 19
rect 90 3 92 7
rect 97 3 99 7
rect 118 3 120 7
rect 128 3 130 7
rect 138 3 140 7
rect 156 5 158 10
rect 163 5 165 10
rect 262 32 264 35
rect 275 32 277 45
rect 295 35 297 53
rect 305 44 307 53
rect 301 42 307 44
rect 301 40 303 42
rect 305 40 307 42
rect 301 38 307 40
rect 312 40 314 53
rect 322 50 324 53
rect 318 48 324 50
rect 318 46 320 48
rect 322 46 324 48
rect 318 44 324 46
rect 312 38 324 40
rect 329 39 331 53
rect 359 56 361 61
rect 339 49 341 52
rect 336 47 342 49
rect 336 45 338 47
rect 340 45 342 47
rect 336 43 342 45
rect 359 44 361 47
rect 262 14 264 19
rect 186 3 188 7
rect 207 3 209 7
rect 217 3 219 7
rect 227 3 229 7
rect 245 5 247 10
rect 252 5 254 10
rect 295 24 297 27
rect 288 22 297 24
rect 305 23 307 38
rect 311 32 317 34
rect 311 30 313 32
rect 315 30 317 32
rect 311 28 317 30
rect 312 23 314 28
rect 322 23 324 38
rect 328 37 334 39
rect 328 35 330 37
rect 332 35 334 37
rect 328 33 334 35
rect 329 23 331 33
rect 339 25 341 43
rect 359 42 365 44
rect 359 40 361 42
rect 363 40 365 42
rect 359 38 365 40
rect 359 35 361 38
rect 288 20 290 22
rect 292 20 294 22
rect 288 18 294 20
rect 359 12 361 17
rect 275 3 277 7
rect 305 3 307 7
rect 312 3 314 7
rect 322 3 324 7
rect 329 3 331 7
rect 339 3 341 7
<< ndif >>
rect -308 96 -297 101
rect -308 94 -306 96
rect -304 94 -297 96
rect -308 92 -297 94
rect -295 99 -288 101
rect -295 97 -292 99
rect -290 97 -288 99
rect -295 95 -288 97
rect -295 92 -290 95
rect -284 94 -277 96
rect -284 92 -282 94
rect -280 92 -277 94
rect -284 90 -277 92
rect -282 87 -277 90
rect -275 95 -270 96
rect -275 91 -267 95
rect -275 89 -272 91
rect -270 89 -267 91
rect -275 87 -267 89
rect -265 87 -260 95
rect -258 91 -250 95
rect -258 89 -255 91
rect -253 89 -250 91
rect -258 87 -250 89
rect -248 87 -243 95
rect -241 93 -233 95
rect -241 91 -238 93
rect -236 91 -233 93
rect -241 89 -233 91
rect -231 93 -224 95
rect -198 94 -193 101
rect -231 91 -228 93
rect -226 91 -224 93
rect -231 89 -224 91
rect -220 92 -213 94
rect -220 90 -218 92
rect -216 90 -213 92
rect -241 87 -235 89
rect -220 88 -213 90
rect -218 81 -213 88
rect -211 88 -203 94
rect -211 86 -208 88
rect -206 86 -203 88
rect -211 84 -203 86
rect -201 91 -193 94
rect -201 89 -198 91
rect -196 89 -193 91
rect -201 87 -193 89
rect -191 99 -183 101
rect -191 97 -188 99
rect -186 97 -183 99
rect -191 87 -183 97
rect -181 99 -174 101
rect -181 97 -178 99
rect -176 97 -174 99
rect -181 92 -174 97
rect -168 94 -163 101
rect -181 90 -178 92
rect -176 90 -174 92
rect -181 87 -174 90
rect -170 92 -163 94
rect -170 90 -168 92
rect -166 90 -163 92
rect -170 88 -163 90
rect -201 84 -196 87
rect -211 81 -206 84
rect -168 81 -163 88
rect -161 81 -156 101
rect -154 95 -147 101
rect -154 85 -145 95
rect -154 83 -151 85
rect -149 83 -145 85
rect -154 81 -145 83
rect -143 92 -136 95
rect -109 94 -104 101
rect -143 90 -140 92
rect -138 90 -136 92
rect -143 88 -136 90
rect -131 92 -124 94
rect -131 90 -129 92
rect -127 90 -124 92
rect -131 88 -124 90
rect -143 81 -138 88
rect -129 81 -124 88
rect -122 88 -114 94
rect -122 86 -119 88
rect -117 86 -114 88
rect -122 84 -114 86
rect -112 91 -104 94
rect -112 89 -109 91
rect -107 89 -104 91
rect -112 87 -104 89
rect -102 99 -94 101
rect -102 97 -99 99
rect -97 97 -94 99
rect -102 87 -94 97
rect -92 99 -85 101
rect -92 97 -89 99
rect -87 97 -85 99
rect -92 92 -85 97
rect -79 94 -74 101
rect -92 90 -89 92
rect -87 90 -85 92
rect -92 87 -85 90
rect -81 92 -74 94
rect -81 90 -79 92
rect -77 90 -74 92
rect -81 88 -74 90
rect -112 84 -107 87
rect -122 81 -117 84
rect -79 81 -74 88
rect -72 81 -67 101
rect -65 95 -58 101
rect -42 95 -35 101
rect -33 99 -25 101
rect -33 97 -30 99
rect -28 97 -25 99
rect -33 95 -25 97
rect -23 95 -15 101
rect -65 85 -56 95
rect -65 83 -62 85
rect -60 83 -56 85
rect -65 81 -56 83
rect -54 92 -47 95
rect -54 90 -51 92
rect -49 90 -47 92
rect -54 88 -47 90
rect -42 88 -37 95
rect -21 92 -15 95
rect -13 99 -6 101
rect -13 97 -10 99
rect -8 97 -6 99
rect -13 95 -6 97
rect -13 92 -8 95
rect 72 98 80 100
rect 72 96 74 98
rect 76 96 80 98
rect 72 94 80 96
rect 82 98 90 100
rect 82 96 85 98
rect 87 96 90 98
rect 82 94 90 96
rect 92 98 99 100
rect 92 96 95 98
rect 97 96 99 98
rect 92 94 99 96
rect 295 95 302 97
rect -21 88 -17 92
rect -54 81 -49 88
rect -42 86 -36 88
rect -42 84 -40 86
rect -38 84 -36 86
rect -42 82 -36 84
rect -23 86 -17 88
rect 2 91 9 93
rect 2 89 4 91
rect 6 89 9 91
rect 2 87 9 89
rect 11 91 19 93
rect 11 89 14 91
rect 16 89 19 91
rect 11 87 19 89
rect 21 87 26 93
rect 28 91 36 93
rect 28 89 31 91
rect 33 89 36 91
rect 28 87 36 89
rect 38 87 43 93
rect 45 91 53 93
rect 45 89 48 91
rect 50 89 53 91
rect 45 87 53 89
rect 55 91 62 93
rect 55 89 58 91
rect 60 89 62 91
rect 103 92 110 94
rect 103 90 105 92
rect 107 90 110 92
rect 55 87 62 89
rect 103 88 110 90
rect 112 92 120 94
rect 112 90 115 92
rect 117 90 120 92
rect 112 88 120 90
rect 122 88 127 94
rect 129 92 137 94
rect 129 90 132 92
rect 134 90 137 92
rect 129 88 137 90
rect 139 88 144 94
rect 146 92 154 94
rect 146 90 149 92
rect 151 90 154 92
rect 146 88 154 90
rect 156 92 163 94
rect 156 90 159 92
rect 161 90 163 92
rect 156 88 163 90
rect 167 92 174 94
rect 167 90 169 92
rect 171 90 174 92
rect 167 88 174 90
rect 176 92 184 94
rect 176 90 179 92
rect 181 90 184 92
rect 176 88 184 90
rect 186 88 191 94
rect 193 92 201 94
rect 193 90 196 92
rect 198 90 201 92
rect 193 88 201 90
rect 203 88 208 94
rect 210 92 218 94
rect 210 90 213 92
rect 215 90 218 92
rect 210 88 218 90
rect 220 92 227 94
rect 220 90 223 92
rect 225 90 227 92
rect 220 88 227 90
rect 231 92 238 94
rect 231 90 233 92
rect 235 90 238 92
rect 231 88 238 90
rect 240 92 248 94
rect 240 90 243 92
rect 245 90 248 92
rect 240 88 248 90
rect 250 88 255 94
rect 257 92 265 94
rect 257 90 260 92
rect 262 90 265 92
rect 257 88 265 90
rect 267 88 272 94
rect 274 92 282 94
rect 274 90 277 92
rect 279 90 282 92
rect 274 88 282 90
rect 284 92 291 94
rect 284 90 287 92
rect 289 90 291 92
rect 295 93 297 95
rect 299 93 302 95
rect 295 91 302 93
rect 304 95 312 97
rect 304 93 307 95
rect 309 93 312 95
rect 304 91 312 93
rect 314 95 322 97
rect 314 93 317 95
rect 319 93 322 95
rect 314 91 322 93
rect 324 95 331 97
rect 324 93 327 95
rect 329 93 331 95
rect 324 91 331 93
rect 336 95 343 97
rect 336 93 338 95
rect 340 93 343 95
rect 336 91 343 93
rect 345 94 353 97
rect 345 91 355 94
rect 284 88 291 90
rect -23 84 -21 86
rect -19 84 -17 86
rect -23 82 -17 84
rect 347 85 355 91
rect 357 85 362 94
rect 364 92 371 94
rect 364 90 367 92
rect 369 90 371 92
rect 364 88 371 90
rect 364 85 369 88
rect 347 83 353 85
rect 347 81 349 83
rect 351 81 353 83
rect 347 79 353 81
rect -289 67 -283 69
rect -289 65 -287 67
rect -285 65 -283 67
rect -289 63 -283 65
rect -305 60 -300 63
rect -307 58 -300 60
rect -307 56 -305 58
rect -303 56 -300 58
rect -307 54 -300 56
rect -298 54 -293 63
rect -291 57 -283 63
rect 81 64 87 66
rect 81 62 83 64
rect 85 62 87 64
rect -227 58 -220 60
rect -291 54 -281 57
rect -289 51 -281 54
rect -279 55 -272 57
rect -279 53 -276 55
rect -274 53 -272 55
rect -279 51 -272 53
rect -267 55 -260 57
rect -267 53 -265 55
rect -263 53 -260 55
rect -267 51 -260 53
rect -258 55 -250 57
rect -258 53 -255 55
rect -253 53 -250 55
rect -258 51 -250 53
rect -248 55 -240 57
rect -248 53 -245 55
rect -243 53 -240 55
rect -248 51 -240 53
rect -238 55 -231 57
rect -238 53 -235 55
rect -233 53 -231 55
rect -227 56 -225 58
rect -223 56 -220 58
rect -227 54 -220 56
rect -218 58 -210 60
rect -218 56 -215 58
rect -213 56 -210 58
rect -218 54 -210 56
rect -208 54 -203 60
rect -201 58 -193 60
rect -201 56 -198 58
rect -196 56 -193 58
rect -201 54 -193 56
rect -191 54 -186 60
rect -184 58 -176 60
rect -184 56 -181 58
rect -179 56 -176 58
rect -184 54 -176 56
rect -174 58 -167 60
rect -174 56 -171 58
rect -169 56 -167 58
rect -174 54 -167 56
rect -163 58 -156 60
rect -163 56 -161 58
rect -159 56 -156 58
rect -163 54 -156 56
rect -154 58 -146 60
rect -154 56 -151 58
rect -149 56 -146 58
rect -154 54 -146 56
rect -144 54 -139 60
rect -137 58 -129 60
rect -137 56 -134 58
rect -132 56 -129 58
rect -137 54 -129 56
rect -127 54 -122 60
rect -120 58 -112 60
rect -120 56 -117 58
rect -115 56 -112 58
rect -120 54 -112 56
rect -110 58 -103 60
rect -110 56 -107 58
rect -105 56 -103 58
rect -110 54 -103 56
rect -99 58 -92 60
rect -99 56 -97 58
rect -95 56 -92 58
rect -99 54 -92 56
rect -90 58 -82 60
rect -90 56 -87 58
rect -85 56 -82 58
rect -90 54 -82 56
rect -80 54 -75 60
rect -73 58 -65 60
rect -73 56 -70 58
rect -68 56 -65 58
rect -73 54 -65 56
rect -63 54 -58 60
rect -56 58 -48 60
rect -56 56 -53 58
rect -51 56 -48 58
rect -56 54 -48 56
rect -46 58 -39 60
rect 2 59 9 61
rect -46 56 -43 58
rect -41 56 -39 58
rect -46 54 -39 56
rect 2 57 4 59
rect 6 57 9 59
rect 2 55 9 57
rect 11 59 19 61
rect 11 57 14 59
rect 16 57 19 59
rect 11 55 19 57
rect 21 55 26 61
rect 28 59 36 61
rect 28 57 31 59
rect 33 57 36 59
rect 28 55 36 57
rect 38 55 43 61
rect 45 59 53 61
rect 45 57 48 59
rect 50 57 53 59
rect 45 55 53 57
rect 55 59 62 61
rect 55 57 58 59
rect 60 57 62 59
rect 55 55 62 57
rect 81 60 87 62
rect 100 64 106 66
rect 100 62 102 64
rect 104 62 106 64
rect 100 60 106 62
rect 113 60 118 67
rect 81 56 85 60
rect -238 51 -231 53
rect -35 52 -28 54
rect -35 50 -33 52
rect -31 50 -28 52
rect -35 48 -28 50
rect -26 52 -18 54
rect -26 50 -23 52
rect -21 50 -18 52
rect -26 48 -18 50
rect -16 52 -8 54
rect -16 50 -12 52
rect -10 50 -8 52
rect -16 48 -8 50
rect 72 53 77 56
rect 70 51 77 53
rect 70 49 72 51
rect 74 49 77 51
rect 70 47 77 49
rect 79 53 85 56
rect 101 53 106 60
rect 111 58 118 60
rect 111 56 113 58
rect 115 56 118 58
rect 111 53 118 56
rect 120 65 129 67
rect 120 63 124 65
rect 126 63 129 65
rect 120 53 129 63
rect 79 47 87 53
rect 89 51 97 53
rect 89 49 92 51
rect 94 49 97 51
rect 89 47 97 49
rect 99 47 106 53
rect 122 47 129 53
rect 131 47 136 67
rect 138 60 143 67
rect 181 64 186 67
rect 171 61 176 64
rect 138 58 145 60
rect 138 56 141 58
rect 143 56 145 58
rect 138 54 145 56
rect 149 58 156 61
rect 149 56 151 58
rect 153 56 156 58
rect 138 47 143 54
rect 149 51 156 56
rect 149 49 151 51
rect 153 49 156 51
rect 149 47 156 49
rect 158 51 166 61
rect 158 49 161 51
rect 163 49 166 51
rect 158 47 166 49
rect 168 59 176 61
rect 168 57 171 59
rect 173 57 176 59
rect 168 54 176 57
rect 178 62 186 64
rect 178 60 181 62
rect 183 60 186 62
rect 178 54 186 60
rect 188 60 193 67
rect 202 60 207 67
rect 188 58 195 60
rect 188 56 191 58
rect 193 56 195 58
rect 188 54 195 56
rect 200 58 207 60
rect 200 56 202 58
rect 204 56 207 58
rect 168 47 173 54
rect 200 53 207 56
rect 209 65 218 67
rect 209 63 213 65
rect 215 63 218 65
rect 209 53 218 63
rect 211 47 218 53
rect 220 47 225 67
rect 227 60 232 67
rect 270 64 275 67
rect 260 61 265 64
rect 227 58 234 60
rect 227 56 230 58
rect 232 56 234 58
rect 227 54 234 56
rect 238 58 245 61
rect 238 56 240 58
rect 242 56 245 58
rect 227 47 232 54
rect 238 51 245 56
rect 238 49 240 51
rect 242 49 245 51
rect 238 47 245 49
rect 247 51 255 61
rect 247 49 250 51
rect 252 49 255 51
rect 247 47 255 49
rect 257 59 265 61
rect 257 57 260 59
rect 262 57 265 59
rect 257 54 265 57
rect 267 62 275 64
rect 267 60 270 62
rect 272 60 275 62
rect 267 54 275 60
rect 277 60 282 67
rect 277 58 284 60
rect 299 59 305 61
rect 277 56 280 58
rect 282 56 284 58
rect 277 54 284 56
rect 288 57 295 59
rect 288 55 290 57
rect 292 55 295 57
rect 257 47 262 54
rect 288 53 295 55
rect 297 57 305 59
rect 297 55 300 57
rect 302 55 305 57
rect 297 53 305 55
rect 307 53 312 61
rect 314 59 322 61
rect 314 57 317 59
rect 319 57 322 59
rect 314 53 322 57
rect 324 53 329 61
rect 331 59 339 61
rect 331 57 334 59
rect 336 57 339 59
rect 331 53 339 57
rect 334 52 339 53
rect 341 58 346 61
rect 341 56 348 58
rect 341 54 344 56
rect 346 54 348 56
rect 341 52 348 54
rect 354 53 359 56
rect 352 51 359 53
rect 352 49 354 51
rect 356 49 359 51
rect 352 47 359 49
rect 361 54 372 56
rect 361 52 368 54
rect 370 52 372 54
rect 361 47 372 52
<< pdif >>
rect -306 132 -299 134
rect -306 130 -303 132
rect -301 131 -299 132
rect -282 134 -277 141
rect -284 132 -277 134
rect -301 130 -297 131
rect -306 113 -297 130
rect -295 126 -290 131
rect -284 130 -282 132
rect -280 130 -277 132
rect -284 128 -277 130
rect -295 124 -288 126
rect -295 122 -292 124
rect -290 122 -288 124
rect -282 123 -277 128
rect -275 139 -267 141
rect -275 137 -272 139
rect -270 137 -267 139
rect -275 125 -267 137
rect -265 125 -260 141
rect -258 129 -250 141
rect -258 127 -255 129
rect -253 127 -250 129
rect -258 125 -250 127
rect -248 125 -243 141
rect -241 139 -234 141
rect -241 137 -238 139
rect -236 137 -234 139
rect -241 129 -234 137
rect -241 125 -235 129
rect -218 129 -213 141
rect -275 123 -270 125
rect -295 117 -288 122
rect -295 115 -292 117
rect -290 115 -288 117
rect -295 113 -288 115
rect -239 121 -235 125
rect -220 127 -213 129
rect -220 125 -218 127
rect -216 125 -213 127
rect -239 113 -233 121
rect -231 119 -226 121
rect -220 120 -213 125
rect -231 117 -224 119
rect -231 115 -228 117
rect -226 115 -224 117
rect -220 118 -218 120
rect -216 118 -213 120
rect -220 116 -213 118
rect -211 139 -202 141
rect -211 137 -207 139
rect -205 137 -202 139
rect -179 139 -165 141
rect -179 138 -172 139
rect -211 129 -202 137
rect -195 129 -190 138
rect -211 116 -200 129
rect -198 120 -190 129
rect -198 118 -195 120
rect -193 118 -190 120
rect -198 116 -190 118
rect -231 113 -224 115
rect -195 113 -190 116
rect -188 113 -183 138
rect -181 137 -172 138
rect -170 137 -165 139
rect -181 132 -165 137
rect -181 130 -172 132
rect -170 130 -165 132
rect -181 113 -165 130
rect -163 131 -155 141
rect -163 129 -160 131
rect -158 129 -155 131
rect -163 124 -155 129
rect -163 122 -160 124
rect -158 122 -155 124
rect -163 113 -155 122
rect -153 139 -145 141
rect -153 137 -150 139
rect -148 137 -145 139
rect -153 132 -145 137
rect -153 130 -150 132
rect -148 130 -145 132
rect -153 113 -145 130
rect -143 126 -138 141
rect -129 129 -124 141
rect -131 127 -124 129
rect -143 124 -136 126
rect -143 122 -140 124
rect -138 122 -136 124
rect -143 117 -136 122
rect -143 115 -140 117
rect -138 115 -136 117
rect -131 125 -129 127
rect -127 125 -124 127
rect -131 120 -124 125
rect -131 118 -129 120
rect -127 118 -124 120
rect -131 116 -124 118
rect -122 139 -113 141
rect -122 137 -118 139
rect -116 137 -113 139
rect -90 139 -76 141
rect -90 138 -83 139
rect -122 129 -113 137
rect -106 129 -101 138
rect -122 116 -111 129
rect -109 120 -101 129
rect -109 118 -106 120
rect -104 118 -101 120
rect -109 116 -101 118
rect -143 113 -136 115
rect -106 113 -101 116
rect -99 113 -94 138
rect -92 137 -83 138
rect -81 137 -76 139
rect -92 132 -76 137
rect -92 130 -83 132
rect -81 130 -76 132
rect -92 113 -76 130
rect -74 131 -66 141
rect -74 129 -71 131
rect -69 129 -66 131
rect -74 124 -66 129
rect -74 122 -71 124
rect -69 122 -66 124
rect -74 113 -66 122
rect -64 139 -56 141
rect -64 137 -61 139
rect -59 137 -56 139
rect -64 132 -56 137
rect -64 130 -61 132
rect -59 130 -56 132
rect -64 113 -56 130
rect -54 126 -49 141
rect -40 134 -35 141
rect -42 132 -35 134
rect -42 130 -40 132
rect -38 130 -35 132
rect -42 128 -35 130
rect -54 124 -47 126
rect -54 122 -51 124
rect -49 122 -47 124
rect -54 117 -47 122
rect -40 120 -35 128
rect -33 120 -28 141
rect -26 139 -17 141
rect -26 137 -21 139
rect -19 137 -17 139
rect -26 131 -17 137
rect 77 135 82 141
rect 75 133 82 135
rect -26 120 -15 131
rect -54 115 -51 117
rect -49 115 -47 117
rect -54 113 -47 115
rect -23 113 -15 120
rect -13 129 -6 131
rect -13 127 -10 129
rect -8 127 -6 129
rect 4 127 9 133
rect -13 122 -6 127
rect -13 120 -10 122
rect -8 120 -6 122
rect 2 125 9 127
rect 2 123 4 125
rect 6 123 9 125
rect 2 121 9 123
rect 11 131 19 133
rect 11 129 14 131
rect 16 129 19 131
rect 11 121 19 129
rect 21 121 26 133
rect 28 125 36 133
rect 28 123 31 125
rect 33 123 36 125
rect 28 121 36 123
rect 38 121 43 133
rect 45 131 52 133
rect 45 129 48 131
rect 50 129 52 131
rect 75 131 77 133
rect 79 131 82 133
rect 75 129 82 131
rect 45 127 52 129
rect 45 121 51 127
rect -13 118 -6 120
rect -13 113 -8 118
rect 47 119 51 121
rect 77 121 82 129
rect 84 121 89 141
rect 91 139 100 141
rect 306 140 315 142
rect 91 137 96 139
rect 98 137 100 139
rect 91 132 100 137
rect 306 138 309 140
rect 311 138 315 140
rect 91 130 96 132
rect 98 130 100 132
rect 91 127 100 130
rect 113 132 120 134
rect 113 130 115 132
rect 117 130 120 132
rect 113 128 120 130
rect 91 121 99 127
rect 47 113 53 119
rect 55 117 62 119
rect 55 115 58 117
rect 60 115 62 117
rect 55 113 62 115
rect 114 122 120 128
rect 122 122 127 134
rect 129 126 137 134
rect 129 124 132 126
rect 134 124 137 126
rect 129 122 137 124
rect 139 122 144 134
rect 146 132 154 134
rect 146 130 149 132
rect 151 130 154 132
rect 146 122 154 130
rect 156 128 161 134
rect 169 128 174 134
rect 156 126 163 128
rect 156 124 159 126
rect 161 124 163 126
rect 156 122 163 124
rect 167 126 174 128
rect 167 124 169 126
rect 171 124 174 126
rect 167 122 174 124
rect 176 132 184 134
rect 176 130 179 132
rect 181 130 184 132
rect 176 122 184 130
rect 186 122 191 134
rect 193 126 201 134
rect 193 124 196 126
rect 198 124 201 126
rect 193 122 201 124
rect 203 122 208 134
rect 210 132 217 134
rect 210 130 213 132
rect 215 130 217 132
rect 210 128 217 130
rect 210 122 216 128
rect 233 128 238 134
rect 114 120 118 122
rect 103 118 110 120
rect 103 116 105 118
rect 107 116 110 118
rect 103 114 110 116
rect 112 114 118 120
rect 212 120 216 122
rect 231 126 238 128
rect 231 124 233 126
rect 235 124 238 126
rect 231 122 238 124
rect 240 132 248 134
rect 240 130 243 132
rect 245 130 248 132
rect 240 122 248 130
rect 250 122 255 134
rect 257 126 265 134
rect 257 124 260 126
rect 262 124 265 126
rect 257 122 265 124
rect 267 122 272 134
rect 274 132 281 134
rect 306 133 315 138
rect 274 130 277 132
rect 279 130 281 132
rect 274 128 281 130
rect 295 131 302 133
rect 295 129 297 131
rect 299 129 302 131
rect 274 122 280 128
rect 295 127 302 129
rect 212 114 218 120
rect 220 118 227 120
rect 220 116 223 118
rect 225 116 227 118
rect 220 114 227 116
rect 276 120 280 122
rect 297 121 302 127
rect 304 124 315 133
rect 317 124 322 142
rect 324 135 329 142
rect 324 133 331 135
rect 324 131 327 133
rect 329 131 331 133
rect 324 129 331 131
rect 324 124 329 129
rect 304 121 312 124
rect 276 114 282 120
rect 284 118 291 120
rect 284 116 287 118
rect 289 116 291 118
rect 284 114 291 116
rect 338 120 343 126
rect 336 118 343 120
rect 336 116 338 118
rect 340 116 343 118
rect 336 114 343 116
rect 345 124 351 126
rect 345 118 353 124
rect 345 116 348 118
rect 350 116 353 118
rect 345 114 353 116
rect 355 118 363 124
rect 355 116 358 118
rect 360 116 363 118
rect 355 114 363 116
rect 365 122 372 124
rect 365 120 368 122
rect 370 120 372 122
rect 365 114 372 120
rect -308 28 -301 34
rect -308 26 -306 28
rect -304 26 -301 28
rect -308 24 -301 26
rect -299 32 -291 34
rect -299 30 -296 32
rect -294 30 -291 32
rect -299 24 -291 30
rect -289 32 -281 34
rect -289 30 -286 32
rect -284 30 -281 32
rect -289 24 -281 30
rect -287 22 -281 24
rect -279 32 -272 34
rect -279 30 -276 32
rect -274 30 -272 32
rect -279 28 -272 30
rect -279 22 -274 28
rect -227 32 -220 34
rect -227 30 -225 32
rect -223 30 -220 32
rect -227 28 -220 30
rect -218 28 -212 34
rect -248 24 -240 27
rect -265 19 -260 24
rect -267 17 -260 19
rect -267 15 -265 17
rect -263 15 -260 17
rect -267 13 -260 15
rect -265 6 -260 13
rect -258 6 -253 24
rect -251 15 -240 24
rect -238 21 -233 27
rect -216 26 -212 28
rect -163 32 -156 34
rect -163 30 -161 32
rect -159 30 -156 32
rect -163 28 -156 30
rect -154 28 -148 34
rect -238 19 -231 21
rect -216 20 -210 26
rect -238 17 -235 19
rect -233 17 -231 19
rect -238 15 -231 17
rect -217 18 -210 20
rect -217 16 -215 18
rect -213 16 -210 18
rect -251 10 -242 15
rect -217 14 -210 16
rect -208 14 -203 26
rect -201 24 -193 26
rect -201 22 -198 24
rect -196 22 -193 24
rect -201 14 -193 22
rect -191 14 -186 26
rect -184 18 -176 26
rect -184 16 -181 18
rect -179 16 -176 18
rect -184 14 -176 16
rect -174 24 -167 26
rect -174 22 -171 24
rect -169 22 -167 24
rect -174 20 -167 22
rect -152 26 -148 28
rect -54 28 -48 34
rect -46 32 -39 34
rect -46 30 -43 32
rect -41 30 -39 32
rect -46 28 -39 30
rect -54 26 -50 28
rect -174 14 -169 20
rect -152 20 -146 26
rect -153 18 -146 20
rect -153 16 -151 18
rect -149 16 -146 18
rect -153 14 -146 16
rect -144 14 -139 26
rect -137 24 -129 26
rect -137 22 -134 24
rect -132 22 -129 24
rect -137 14 -129 22
rect -127 14 -122 26
rect -120 18 -112 26
rect -120 16 -117 18
rect -115 16 -112 18
rect -120 14 -112 16
rect -110 24 -103 26
rect -110 22 -107 24
rect -105 22 -103 24
rect -110 20 -103 22
rect -99 24 -92 26
rect -99 22 -97 24
rect -95 22 -92 24
rect -99 20 -92 22
rect -110 14 -105 20
rect -97 14 -92 20
rect -90 18 -82 26
rect -90 16 -87 18
rect -85 16 -82 18
rect -90 14 -82 16
rect -80 14 -75 26
rect -73 24 -65 26
rect -73 22 -70 24
rect -68 22 -65 24
rect -73 14 -65 22
rect -63 14 -58 26
rect -56 20 -50 26
rect 2 33 9 35
rect 2 31 4 33
rect 6 31 9 33
rect 2 29 9 31
rect 11 29 17 35
rect -35 21 -27 27
rect -56 18 -49 20
rect -56 16 -53 18
rect -51 16 -49 18
rect -56 14 -49 16
rect -36 18 -27 21
rect -36 16 -34 18
rect -32 16 -27 18
rect -251 8 -247 10
rect -245 8 -242 10
rect -36 11 -27 16
rect -36 9 -34 11
rect -32 9 -27 11
rect -251 6 -242 8
rect -36 7 -27 9
rect -25 7 -20 27
rect -18 19 -13 27
rect 13 27 17 29
rect 72 30 77 35
rect 70 28 77 30
rect 13 21 19 27
rect 12 19 19 21
rect -18 17 -11 19
rect -18 15 -15 17
rect -13 15 -11 17
rect 12 17 14 19
rect 16 17 19 19
rect 12 15 19 17
rect 21 15 26 27
rect 28 25 36 27
rect 28 23 31 25
rect 33 23 36 25
rect 28 15 36 23
rect 38 15 43 27
rect 45 19 53 27
rect 45 17 48 19
rect 50 17 53 19
rect 45 15 53 17
rect 55 25 62 27
rect 55 23 58 25
rect 60 23 62 25
rect 55 21 62 23
rect 70 26 72 28
rect 74 26 77 28
rect 70 21 77 26
rect 55 15 60 21
rect 70 19 72 21
rect 74 19 77 21
rect 70 17 77 19
rect 79 28 87 35
rect 111 33 118 35
rect 111 31 113 33
rect 115 31 118 33
rect 79 17 90 28
rect -18 13 -11 15
rect -18 7 -13 13
rect 81 11 90 17
rect 81 9 83 11
rect 85 9 90 11
rect 81 7 90 9
rect 92 7 97 28
rect 99 20 104 28
rect 111 26 118 31
rect 111 24 113 26
rect 115 24 118 26
rect 111 22 118 24
rect 99 18 106 20
rect 99 16 102 18
rect 104 16 106 18
rect 99 14 106 16
rect 99 7 104 14
rect 113 7 118 22
rect 120 18 128 35
rect 120 16 123 18
rect 125 16 128 18
rect 120 11 128 16
rect 120 9 123 11
rect 125 9 128 11
rect 120 7 128 9
rect 130 26 138 35
rect 130 24 133 26
rect 135 24 138 26
rect 130 19 138 24
rect 130 17 133 19
rect 135 17 138 19
rect 130 7 138 17
rect 140 18 156 35
rect 140 16 145 18
rect 147 16 156 18
rect 140 11 156 16
rect 140 9 145 11
rect 147 10 156 11
rect 158 10 163 35
rect 165 32 170 35
rect 200 33 207 35
rect 165 30 173 32
rect 165 28 168 30
rect 170 28 173 30
rect 165 19 173 28
rect 175 19 186 32
rect 165 10 170 19
rect 177 11 186 19
rect 147 9 154 10
rect 140 7 154 9
rect 177 9 180 11
rect 182 9 186 11
rect 177 7 186 9
rect 188 30 195 32
rect 188 28 191 30
rect 193 28 195 30
rect 188 23 195 28
rect 188 21 191 23
rect 193 21 195 23
rect 200 31 202 33
rect 204 31 207 33
rect 200 26 207 31
rect 200 24 202 26
rect 204 24 207 26
rect 200 22 207 24
rect 188 19 195 21
rect 188 7 193 19
rect 202 7 207 22
rect 209 18 217 35
rect 209 16 212 18
rect 214 16 217 18
rect 209 11 217 16
rect 209 9 212 11
rect 214 9 217 11
rect 209 7 217 9
rect 219 26 227 35
rect 219 24 222 26
rect 224 24 227 26
rect 219 19 227 24
rect 219 17 222 19
rect 224 17 227 19
rect 219 7 227 17
rect 229 18 245 35
rect 229 16 234 18
rect 236 16 245 18
rect 229 11 245 16
rect 229 9 234 11
rect 236 10 245 11
rect 247 10 252 35
rect 254 32 259 35
rect 288 33 295 35
rect 254 30 262 32
rect 254 28 257 30
rect 259 28 262 30
rect 254 19 262 28
rect 264 19 275 32
rect 254 10 259 19
rect 266 11 275 19
rect 236 9 243 10
rect 229 7 243 9
rect 266 9 269 11
rect 271 9 275 11
rect 266 7 275 9
rect 277 30 284 32
rect 277 28 280 30
rect 282 28 284 30
rect 288 31 290 33
rect 292 31 295 33
rect 288 29 295 31
rect 277 23 284 28
rect 290 27 295 29
rect 297 27 303 35
rect 277 21 280 23
rect 282 21 284 23
rect 277 19 284 21
rect 299 23 303 27
rect 352 33 359 35
rect 352 31 354 33
rect 356 31 359 33
rect 352 26 359 31
rect 334 23 339 25
rect 277 7 282 19
rect 299 19 305 23
rect 298 11 305 19
rect 298 9 300 11
rect 302 9 305 11
rect 298 7 305 9
rect 307 7 312 23
rect 314 21 322 23
rect 314 19 317 21
rect 319 19 322 21
rect 314 7 322 19
rect 324 7 329 23
rect 331 11 339 23
rect 331 9 334 11
rect 336 9 339 11
rect 331 7 339 9
rect 341 20 346 25
rect 352 24 354 26
rect 356 24 359 26
rect 352 22 359 24
rect 341 18 348 20
rect 341 16 344 18
rect 346 16 348 18
rect 354 17 359 22
rect 361 18 370 35
rect 361 17 365 18
rect 341 14 348 16
rect 341 7 346 14
rect 363 16 365 17
rect 367 16 370 18
rect 363 14 370 16
<< alu1 >>
rect -312 143 376 147
rect -312 142 106 143
rect -312 140 -305 142
rect -303 140 -293 142
rect -291 140 -11 142
rect -9 140 57 142
rect 59 141 106 142
rect 108 141 222 143
rect 224 141 286 143
rect 288 141 298 143
rect 300 141 339 143
rect 341 141 353 143
rect 355 141 367 143
rect 369 141 376 143
rect 59 140 376 141
rect -312 139 100 140
rect -284 132 -271 133
rect -284 130 -282 132
rect -280 130 -271 132
rect -284 129 -271 130
rect -300 124 -288 126
rect -300 122 -292 124
rect -290 122 -288 124
rect -300 120 -288 122
rect -292 117 -288 120
rect -290 115 -288 117
rect -308 108 -296 110
rect -308 106 -306 108
rect -304 106 -299 108
rect -297 106 -296 108
rect -308 104 -296 106
rect -300 96 -296 104
rect -292 103 -288 115
rect -292 101 -291 103
rect -289 101 -288 103
rect -292 99 -288 101
rect -290 97 -288 99
rect -292 88 -288 97
rect -284 108 -280 129
rect -229 128 -224 134
rect -229 126 -228 128
rect -226 126 -224 128
rect -284 106 -283 108
rect -281 106 -280 108
rect -284 96 -280 106
rect -229 125 -224 126
rect -237 121 -224 125
rect -220 129 -207 133
rect -131 129 -118 133
rect -10 133 -6 134
rect -19 129 -6 133
rect -220 127 -215 129
rect -220 125 -218 127
rect -216 125 -215 127
rect -131 127 -126 129
rect -220 120 -215 125
rect -220 118 -218 120
rect -216 118 -215 120
rect -268 116 -256 118
rect -268 114 -263 116
rect -261 114 -256 116
rect -268 113 -256 114
rect -266 112 -256 113
rect -266 111 -264 112
rect -268 104 -264 111
rect -244 108 -238 110
rect -244 106 -241 108
rect -239 106 -238 108
rect -244 101 -238 106
rect -244 100 -231 101
rect -244 98 -243 100
rect -241 98 -231 100
rect -244 97 -231 98
rect -284 94 -279 96
rect -284 92 -282 94
rect -280 92 -279 94
rect -284 90 -279 92
rect -284 88 -280 90
rect -220 116 -215 118
rect -220 96 -216 116
rect -189 116 -151 117
rect -189 114 -160 116
rect -158 114 -151 116
rect -189 113 -151 114
rect -189 110 -184 113
rect -192 108 -184 110
rect -192 106 -191 108
rect -189 106 -184 108
rect -192 104 -184 106
rect -174 108 -159 109
rect -174 106 -172 108
rect -170 106 -165 108
rect -163 106 -159 108
rect -174 105 -159 106
rect -220 94 -219 96
rect -217 94 -216 96
rect -220 92 -215 94
rect -172 99 -168 105
rect -141 124 -135 126
rect -141 122 -140 124
rect -138 122 -135 124
rect -141 117 -135 122
rect -141 115 -140 117
rect -138 115 -135 117
rect -141 113 -135 115
rect -172 97 -171 99
rect -169 97 -168 99
rect -172 96 -168 97
rect -139 99 -135 113
rect -139 97 -138 99
rect -136 97 -135 99
rect -139 93 -135 97
rect -220 90 -218 92
rect -216 90 -215 92
rect -220 88 -215 90
rect -157 92 -135 93
rect -157 90 -140 92
rect -138 90 -135 92
rect -157 89 -135 90
rect -131 125 -129 127
rect -127 125 -126 127
rect -131 120 -126 125
rect -131 118 -129 120
rect -127 118 -126 120
rect -131 116 -126 118
rect -131 114 -130 116
rect -128 114 -127 116
rect -131 94 -127 114
rect -100 113 -62 117
rect -100 110 -95 113
rect -103 108 -95 110
rect -103 106 -102 108
rect -100 106 -98 108
rect -96 106 -95 108
rect -103 104 -95 106
rect -85 108 -70 109
rect -85 106 -83 108
rect -81 106 -76 108
rect -74 106 -70 108
rect -85 105 -70 106
rect -131 92 -126 94
rect -83 96 -79 105
rect -52 124 -46 126
rect -52 122 -51 124
rect -49 123 -46 124
rect -42 123 -38 126
rect -49 122 -38 123
rect -52 119 -38 122
rect -52 117 -46 119
rect -52 115 -51 117
rect -49 115 -46 117
rect -52 113 -46 115
rect -42 117 -38 119
rect -42 115 -21 117
rect -42 113 -37 115
rect -35 113 -21 115
rect -50 93 -46 113
rect -42 108 -21 109
rect -42 106 -27 108
rect -25 106 -21 108
rect -42 105 -21 106
rect -8 127 -6 129
rect 57 132 62 134
rect 57 130 58 132
rect 60 130 62 132
rect -10 122 -6 127
rect 57 126 62 130
rect -8 120 -6 122
rect -42 99 -38 105
rect -10 110 -6 120
rect -10 108 -9 110
rect -7 108 -6 110
rect -10 101 -6 108
rect -42 97 -41 99
rect -39 97 -38 99
rect -42 96 -38 97
rect -11 99 -6 101
rect -11 97 -10 99
rect -8 97 -6 99
rect -11 95 -6 97
rect 2 125 8 126
rect 57 125 58 126
rect 2 123 4 125
rect 6 123 15 125
rect 2 121 15 123
rect 49 124 58 125
rect 60 124 62 126
rect 49 121 62 124
rect 72 133 81 134
rect 72 131 77 133
rect 79 131 81 133
rect 72 130 81 131
rect -131 90 -129 92
rect -127 90 -126 92
rect -131 88 -126 90
rect -68 92 -46 93
rect -68 90 -51 92
rect -49 90 -46 92
rect -68 89 -46 90
rect 2 92 6 121
rect 25 111 31 117
rect 16 110 31 111
rect 16 108 18 110
rect 20 108 27 110
rect 29 108 31 110
rect 16 105 31 108
rect 42 108 48 110
rect 42 106 45 108
rect 47 106 48 108
rect 42 102 48 106
rect 42 99 54 102
rect 42 97 48 99
rect 50 97 54 99
rect 42 96 54 97
rect 2 91 8 92
rect 2 89 4 91
rect 6 89 8 91
rect 2 88 8 89
rect 72 113 76 130
rect 103 132 108 134
rect 103 130 104 132
rect 106 130 108 132
rect 103 127 108 130
rect 222 131 227 135
rect 222 129 224 131
rect 226 129 227 131
rect 291 139 295 140
rect 286 132 291 135
rect 286 130 288 132
rect 290 130 291 132
rect 222 127 227 129
rect 286 127 291 130
rect 88 125 92 126
rect 88 123 89 125
rect 91 123 92 125
rect 88 121 92 123
rect 103 125 105 127
rect 107 126 108 127
rect 157 126 163 127
rect 107 125 116 126
rect 103 122 116 125
rect 150 124 159 126
rect 161 124 163 126
rect 150 122 163 124
rect 72 111 73 113
rect 75 111 76 113
rect 80 117 92 121
rect 96 117 100 118
rect 80 116 84 117
rect 80 114 81 116
rect 83 114 84 116
rect 80 112 84 114
rect 96 115 97 117
rect 99 115 100 117
rect 72 108 76 111
rect 96 110 100 115
rect 72 104 84 108
rect 88 107 100 110
rect 88 105 91 107
rect 93 105 100 107
rect 88 104 100 105
rect 80 99 84 104
rect 80 98 89 99
rect 80 96 85 98
rect 87 96 89 98
rect 80 95 89 96
rect 117 109 123 111
rect 117 107 118 109
rect 120 107 123 109
rect 117 103 123 107
rect 111 101 123 103
rect 111 99 117 101
rect 119 99 123 101
rect 111 97 123 99
rect 134 112 140 118
rect 134 111 149 112
rect 134 110 145 111
rect 134 108 140 110
rect 142 109 145 110
rect 147 109 149 111
rect 142 108 149 109
rect 134 106 149 108
rect 159 110 163 122
rect 159 108 160 110
rect 162 108 163 110
rect 159 93 163 108
rect 157 92 163 93
rect 157 90 159 92
rect 161 90 163 92
rect 157 89 163 90
rect 167 126 173 127
rect 222 126 223 127
rect 167 124 169 126
rect 171 124 180 126
rect 167 122 180 124
rect 214 125 223 126
rect 225 125 227 127
rect 214 122 227 125
rect 231 126 237 127
rect 286 126 287 127
rect 231 124 233 126
rect 235 124 244 126
rect 231 122 244 124
rect 278 125 287 126
rect 289 125 291 127
rect 278 122 291 125
rect 295 131 308 134
rect 295 129 297 131
rect 299 130 308 131
rect 167 93 171 122
rect 190 112 196 118
rect 181 111 196 112
rect 181 109 183 111
rect 185 110 196 111
rect 185 109 188 110
rect 181 108 188 109
rect 190 108 196 110
rect 181 106 196 108
rect 207 109 213 111
rect 207 107 210 109
rect 212 107 213 109
rect 207 103 213 107
rect 207 101 219 103
rect 207 99 212 101
rect 214 99 219 101
rect 207 97 219 99
rect 167 92 173 93
rect 167 90 169 92
rect 171 90 173 92
rect 167 89 173 90
rect 231 101 235 122
rect 231 99 232 101
rect 234 99 235 101
rect 231 93 235 99
rect 254 113 260 118
rect 254 112 257 113
rect 245 111 257 112
rect 259 111 260 113
rect 245 109 247 111
rect 249 109 260 111
rect 245 106 260 109
rect 271 109 277 111
rect 271 107 274 109
rect 276 107 277 109
rect 271 103 277 107
rect 271 100 283 103
rect 271 98 280 100
rect 282 98 283 100
rect 271 97 283 98
rect 231 92 237 93
rect 231 90 233 92
rect 235 90 237 92
rect 231 89 237 90
rect 295 113 299 129
rect 295 111 296 113
rect 298 111 299 113
rect 295 97 299 111
rect 319 126 323 127
rect 319 124 320 126
rect 322 124 323 126
rect 319 118 323 124
rect 310 117 323 118
rect 310 115 314 117
rect 316 115 323 117
rect 310 114 323 115
rect 327 110 331 119
rect 318 109 331 110
rect 318 107 324 109
rect 326 107 328 109
rect 330 107 331 109
rect 318 106 331 107
rect 327 105 331 106
rect 336 118 340 127
rect 336 116 338 118
rect 295 95 300 97
rect 295 93 297 95
rect 299 93 300 95
rect 295 89 300 93
rect 336 100 340 116
rect 351 133 364 135
rect 351 131 355 133
rect 357 131 364 133
rect 351 129 364 131
rect 351 126 357 129
rect 351 124 353 126
rect 355 124 357 126
rect 351 122 357 124
rect 368 109 372 111
rect 368 107 369 109
rect 371 107 372 109
rect 336 98 337 100
rect 339 98 340 100
rect 336 95 340 98
rect 336 93 338 95
rect 340 93 348 95
rect 336 89 348 93
rect 368 102 372 107
rect 359 101 372 102
rect 359 99 364 101
rect 366 99 372 101
rect 359 97 372 99
rect 70 83 376 84
rect -312 82 298 83
rect -312 80 -305 82
rect -303 80 -293 82
rect -291 80 -11 82
rect -9 80 75 82
rect 77 80 95 82
rect 97 81 298 82
rect 300 81 326 83
rect 328 81 339 83
rect 341 81 349 83
rect 351 81 376 83
rect 97 80 376 81
rect -312 68 376 80
rect -312 67 -33 68
rect -312 65 -287 67
rect -285 65 -277 67
rect -275 65 -264 67
rect -262 65 -236 67
rect -234 66 -33 67
rect -31 66 -13 68
rect -11 66 73 68
rect 75 66 355 68
rect 357 66 367 68
rect 369 66 376 68
rect -234 65 376 66
rect -312 64 -7 65
rect -308 49 -295 51
rect -308 47 -302 49
rect -300 47 -295 49
rect -308 46 -295 47
rect -308 41 -304 46
rect -284 55 -272 59
rect -284 53 -276 55
rect -274 53 -272 55
rect -276 50 -272 53
rect -276 48 -275 50
rect -273 48 -272 50
rect -308 39 -307 41
rect -305 39 -304 41
rect -308 37 -304 39
rect -293 24 -287 26
rect -293 22 -291 24
rect -289 22 -287 24
rect -293 19 -287 22
rect -300 17 -287 19
rect -300 15 -293 17
rect -291 15 -287 17
rect -300 13 -287 15
rect -276 32 -272 48
rect -236 55 -231 59
rect -236 53 -235 55
rect -233 53 -231 55
rect -236 51 -231 53
rect -274 30 -272 32
rect -276 21 -272 30
rect -267 42 -263 43
rect -267 41 -254 42
rect -267 39 -266 41
rect -264 39 -262 41
rect -260 39 -254 41
rect -267 38 -254 39
rect -267 29 -263 38
rect -259 33 -246 34
rect -259 31 -252 33
rect -250 31 -246 33
rect -259 30 -246 31
rect -259 24 -255 30
rect -259 22 -258 24
rect -256 22 -255 24
rect -259 21 -255 22
rect -235 37 -231 51
rect -235 35 -234 37
rect -232 35 -231 37
rect -235 19 -231 35
rect -173 58 -167 59
rect -173 56 -171 58
rect -169 56 -167 58
rect -173 55 -167 56
rect -219 50 -207 51
rect -219 48 -218 50
rect -216 48 -207 50
rect -219 45 -207 48
rect -213 41 -207 45
rect -213 39 -212 41
rect -210 39 -207 41
rect -213 37 -207 39
rect -196 39 -181 42
rect -196 37 -185 39
rect -183 37 -181 39
rect -196 35 -195 37
rect -193 36 -181 37
rect -193 35 -190 36
rect -196 30 -190 35
rect -171 49 -167 55
rect -171 47 -170 49
rect -168 47 -167 49
rect -171 26 -167 47
rect -109 58 -103 59
rect -109 56 -107 58
rect -105 56 -103 58
rect -109 55 -103 56
rect -155 49 -143 51
rect -155 47 -150 49
rect -148 47 -143 49
rect -155 45 -143 47
rect -149 41 -143 45
rect -149 39 -148 41
rect -146 39 -143 41
rect -149 37 -143 39
rect -132 40 -117 42
rect -132 38 -126 40
rect -124 39 -117 40
rect -124 38 -121 39
rect -132 37 -121 38
rect -119 37 -117 39
rect -132 36 -117 37
rect -132 30 -126 36
rect -107 26 -103 55
rect -244 17 -235 18
rect -233 17 -231 19
rect -244 14 -231 17
rect -227 23 -214 26
rect -227 21 -225 23
rect -223 22 -214 23
rect -180 24 -167 26
rect -180 22 -171 24
rect -169 22 -167 24
rect -223 21 -222 22
rect -173 21 -167 22
rect -163 23 -150 26
rect -163 21 -161 23
rect -159 22 -150 23
rect -116 24 -103 26
rect -116 22 -107 24
rect -105 22 -103 24
rect -159 21 -158 22
rect -109 21 -103 22
rect -99 58 -93 59
rect -99 56 -97 58
rect -95 56 -93 58
rect -99 55 -93 56
rect -99 40 -95 55
rect -99 38 -98 40
rect -96 38 -95 40
rect -99 26 -95 38
rect -85 40 -70 42
rect -85 39 -78 40
rect -85 37 -83 39
rect -81 38 -78 39
rect -76 38 -70 40
rect -81 37 -70 38
rect -85 36 -70 37
rect -76 30 -70 36
rect -59 49 -47 51
rect -59 47 -55 49
rect -53 47 -47 49
rect -59 45 -47 47
rect -59 41 -53 45
rect -59 39 -56 41
rect -54 39 -53 41
rect -59 37 -53 39
rect -25 52 -16 53
rect -25 50 -23 52
rect -21 50 -16 52
rect -25 49 -16 50
rect -20 44 -16 49
rect -36 43 -24 44
rect -36 41 -29 43
rect -27 41 -24 43
rect -36 38 -24 41
rect -20 40 -8 44
rect -36 33 -32 38
rect -12 37 -8 40
rect -36 31 -35 33
rect -33 31 -32 33
rect -20 34 -16 36
rect -20 32 -19 34
rect -17 32 -16 34
rect -20 31 -16 32
rect -36 30 -32 31
rect -28 27 -16 31
rect -12 35 -11 37
rect -9 35 -8 37
rect -99 24 -86 26
rect -99 22 -97 24
rect -95 22 -86 24
rect -52 23 -39 26
rect -52 22 -43 23
rect -99 21 -93 22
rect -44 21 -43 22
rect -41 21 -39 23
rect -28 25 -24 27
rect -28 23 -27 25
rect -25 23 -24 25
rect -28 22 -24 23
rect -227 18 -222 21
rect -163 19 -158 21
rect -227 16 -226 18
rect -224 16 -222 18
rect -227 13 -222 16
rect -231 8 -227 9
rect -163 17 -162 19
rect -160 17 -158 19
rect -163 13 -158 17
rect -44 18 -39 21
rect -44 16 -42 18
rect -40 16 -39 18
rect -44 14 -39 16
rect -12 18 -8 35
rect 56 59 62 60
rect 56 57 58 59
rect 60 57 62 59
rect 56 56 62 57
rect 10 51 22 52
rect 10 49 14 51
rect 16 49 22 51
rect 10 46 22 49
rect 16 42 22 46
rect 16 40 17 42
rect 19 40 22 42
rect 16 38 22 40
rect 33 40 48 43
rect 33 38 35 40
rect 37 38 44 40
rect 46 38 48 40
rect 33 37 48 38
rect 33 31 39 37
rect 58 27 62 56
rect 110 58 132 59
rect 110 56 113 58
rect 115 56 132 58
rect 110 55 132 56
rect 190 58 195 60
rect 190 56 191 58
rect 193 56 195 58
rect -17 17 -8 18
rect -17 15 -15 17
rect -13 15 -8 17
rect -17 14 -8 15
rect 2 24 15 27
rect 2 22 4 24
rect 6 23 15 24
rect 49 25 62 27
rect 49 23 58 25
rect 60 23 62 25
rect 6 22 7 23
rect 56 22 62 23
rect 70 51 75 53
rect 70 49 72 51
rect 74 49 75 51
rect 70 47 75 49
rect 102 51 106 52
rect 102 49 103 51
rect 105 49 106 51
rect 70 40 74 47
rect 70 38 71 40
rect 73 38 74 40
rect 70 28 74 38
rect 102 43 106 49
rect 70 26 72 28
rect 2 18 7 22
rect 70 21 74 26
rect 2 16 4 18
rect 6 16 7 18
rect 2 14 7 16
rect 70 19 72 21
rect 85 42 106 43
rect 85 40 89 42
rect 91 40 106 42
rect 85 39 106 40
rect 110 35 114 55
rect 85 33 99 35
rect 101 33 106 35
rect 85 31 106 33
rect 102 29 106 31
rect 110 33 116 35
rect 110 31 113 33
rect 115 31 116 33
rect 110 29 116 31
rect 102 26 116 29
rect 102 25 113 26
rect 102 22 106 25
rect 110 24 113 25
rect 115 24 116 26
rect 110 22 116 24
rect 143 43 147 52
rect 190 54 195 56
rect 134 42 149 43
rect 134 40 138 42
rect 140 40 145 42
rect 147 40 149 42
rect 134 39 149 40
rect 159 42 167 44
rect 159 40 160 42
rect 162 40 164 42
rect 166 40 167 42
rect 159 38 167 40
rect 159 35 164 38
rect 126 31 164 35
rect 191 34 195 54
rect 191 32 192 34
rect 194 32 195 34
rect 190 30 195 32
rect 190 28 191 30
rect 193 28 195 30
rect 190 23 195 28
rect 190 21 191 23
rect 193 21 195 23
rect 199 58 221 59
rect 199 56 202 58
rect 204 56 221 58
rect 199 55 221 56
rect 279 58 284 60
rect 279 56 280 58
rect 282 56 284 58
rect 199 51 203 55
rect 199 49 200 51
rect 202 49 203 51
rect 199 35 203 49
rect 232 51 236 52
rect 232 49 233 51
rect 235 49 236 51
rect 199 33 205 35
rect 199 31 202 33
rect 204 31 205 33
rect 199 26 205 31
rect 199 24 202 26
rect 204 24 205 26
rect 199 22 205 24
rect 232 43 236 49
rect 279 54 284 56
rect 280 52 281 54
rect 283 52 284 54
rect 223 42 238 43
rect 223 40 227 42
rect 229 40 234 42
rect 236 40 238 42
rect 223 39 238 40
rect 248 42 256 44
rect 248 40 253 42
rect 255 40 256 42
rect 248 38 256 40
rect 248 35 253 38
rect 215 34 253 35
rect 215 32 222 34
rect 224 32 253 34
rect 215 31 253 32
rect 280 32 284 52
rect 279 30 284 32
rect 344 58 348 60
rect 343 56 348 58
rect 343 54 344 56
rect 346 54 348 56
rect 343 52 348 54
rect 295 50 308 51
rect 295 48 305 50
rect 307 48 308 50
rect 295 47 308 48
rect 302 42 308 47
rect 302 40 303 42
rect 305 40 308 42
rect 302 38 308 40
rect 328 37 332 44
rect 328 36 330 37
rect 320 35 330 36
rect 320 34 332 35
rect 320 32 325 34
rect 327 32 332 34
rect 320 30 332 32
rect 279 28 280 30
rect 282 28 284 30
rect 279 23 284 28
rect 190 19 195 21
rect 279 21 280 23
rect 282 21 284 23
rect 279 19 284 21
rect 70 15 83 19
rect 70 14 74 15
rect 182 15 195 19
rect 271 15 284 19
rect 288 23 301 27
rect 288 22 293 23
rect 344 42 348 52
rect 344 40 345 42
rect 347 40 348 42
rect 288 20 290 22
rect 292 20 293 22
rect 288 14 293 20
rect 344 19 348 40
rect 352 51 356 60
rect 352 49 354 51
rect 352 47 356 49
rect 352 45 353 47
rect 355 45 356 47
rect 352 33 356 45
rect 360 44 364 52
rect 360 42 372 44
rect 360 40 361 42
rect 363 40 368 42
rect 370 40 372 42
rect 360 38 372 40
rect 352 31 354 33
rect 352 28 356 31
rect 352 26 364 28
rect 352 24 354 26
rect 356 24 364 26
rect 352 22 364 24
rect 335 18 348 19
rect 335 16 344 18
rect 346 16 348 18
rect 335 15 348 16
rect -36 8 376 9
rect -312 7 5 8
rect -312 5 -305 7
rect -303 5 -291 7
rect -289 5 -277 7
rect -275 5 -236 7
rect -234 5 -224 7
rect -222 5 -160 7
rect -158 5 -44 7
rect -42 6 5 7
rect 7 6 73 8
rect 75 6 355 8
rect 357 6 367 8
rect 369 6 376 8
rect -42 5 376 6
rect -312 1 376 5
<< alu2 >>
rect 212 136 235 140
rect 57 132 62 134
rect 212 133 216 136
rect 57 130 58 132
rect 60 130 62 132
rect -308 116 -260 117
rect -308 114 -263 116
rect -261 114 -260 116
rect -308 113 -260 114
rect -161 116 -127 117
rect -161 114 -160 116
rect -158 114 -130 116
rect -128 114 -127 116
rect -161 113 -127 114
rect -308 108 -303 113
rect -10 110 31 111
rect -308 106 -306 108
rect -304 106 -303 108
rect -308 43 -303 106
rect -284 108 -95 109
rect -284 106 -283 108
rect -281 106 -98 108
rect -96 106 -95 108
rect -10 108 -9 110
rect -7 108 27 110
rect 29 108 31 110
rect -10 107 31 108
rect -284 105 -95 106
rect -292 103 -288 104
rect -292 101 -291 103
rect -289 101 -288 103
rect -292 100 -240 101
rect -292 98 -243 100
rect -241 98 -240 100
rect -292 97 -240 98
rect -172 99 -168 101
rect -172 97 -171 99
rect -169 97 -168 99
rect -220 96 -216 97
rect -220 94 -219 96
rect -217 94 -216 96
rect -220 83 -216 94
rect -172 92 -168 97
rect -139 99 52 100
rect -139 97 -138 99
rect -136 97 -134 99
rect -132 97 -41 99
rect -39 97 48 99
rect 50 97 52 99
rect -139 96 52 97
rect -172 88 -47 92
rect -220 79 -80 83
rect -276 50 -215 51
rect -276 48 -275 50
rect -273 48 -218 50
rect -216 48 -215 50
rect -276 47 -215 48
rect -171 49 -143 51
rect -171 47 -170 49
rect -168 47 -150 49
rect -148 47 -143 49
rect -171 45 -143 47
rect -308 41 -263 43
rect -85 42 -80 79
rect -53 51 -47 88
rect 57 81 62 130
rect 88 132 216 133
rect 231 133 235 136
rect 231 132 291 133
rect 88 130 104 132
rect 106 130 216 132
rect 88 129 216 130
rect 221 131 227 132
rect 221 129 224 131
rect 226 129 227 131
rect 231 130 288 132
rect 290 130 291 132
rect 231 129 291 130
rect 88 125 92 129
rect 221 125 227 129
rect 88 123 89 125
rect 91 123 92 125
rect 88 122 92 123
rect 96 121 227 125
rect 318 126 357 127
rect 318 124 320 126
rect 322 124 353 126
rect 355 124 357 126
rect 318 123 357 124
rect 96 117 100 121
rect 318 118 323 123
rect -12 76 62 81
rect 72 113 76 116
rect 96 115 97 117
rect 99 115 100 117
rect 96 113 100 115
rect 310 117 323 118
rect 310 115 311 117
rect 313 115 323 117
rect 310 114 323 115
rect 255 113 299 114
rect 72 111 73 113
rect 75 111 76 113
rect -59 49 -41 51
rect -59 47 -55 49
rect -53 47 -41 49
rect -59 45 -41 47
rect -308 39 -307 41
rect -305 39 -266 41
rect -264 39 -263 41
rect -308 37 -263 39
rect -132 40 -95 42
rect -132 38 -126 40
rect -124 38 -98 40
rect -96 38 -95 40
rect -235 37 -191 38
rect -235 35 -234 37
rect -232 35 -195 37
rect -193 35 -191 37
rect -132 36 -95 38
rect -85 40 -73 42
rect -85 38 -78 40
rect -76 38 -73 40
rect -85 36 -73 38
rect -12 37 -8 76
rect 72 71 76 111
rect 137 110 149 112
rect 137 108 140 110
rect 142 108 149 110
rect 137 106 149 108
rect 159 110 196 112
rect 255 111 257 113
rect 259 111 296 113
rect 298 111 299 113
rect 255 110 299 111
rect 159 108 160 110
rect 162 108 188 110
rect 190 108 196 110
rect 159 106 196 108
rect 327 109 372 111
rect 327 107 328 109
rect 330 107 369 109
rect 371 107 372 109
rect 105 101 123 103
rect 105 99 117 101
rect 119 99 123 101
rect 105 97 123 99
rect -12 35 -11 37
rect -9 35 -8 37
rect -235 34 -191 35
rect -259 33 -246 34
rect -259 31 -249 33
rect -247 31 -246 33
rect -259 30 -246 31
rect -36 33 -32 35
rect -36 31 -35 33
rect -33 31 -32 33
rect -12 32 -8 35
rect 2 66 76 71
rect -259 25 -254 30
rect -36 27 -32 31
rect -293 24 -254 25
rect -293 22 -291 24
rect -289 22 -258 24
rect -256 22 -254 24
rect -293 21 -254 22
rect -163 23 -32 27
rect -28 25 -24 26
rect -28 23 -27 25
rect -25 23 -24 25
rect -163 19 -157 23
rect -28 19 -24 23
rect -227 18 -167 19
rect -227 16 -226 18
rect -224 16 -167 18
rect -163 17 -162 19
rect -160 17 -157 19
rect -163 16 -157 17
rect -152 18 -24 19
rect -152 16 -42 18
rect -40 16 -24 18
rect -227 15 -167 16
rect -171 12 -167 15
rect -152 15 -24 16
rect 2 18 7 66
rect 111 60 117 97
rect 144 69 149 106
rect 327 105 372 107
rect 207 101 235 103
rect 207 99 212 101
rect 214 99 232 101
rect 234 99 235 101
rect 207 97 235 99
rect 279 100 340 101
rect 279 98 280 100
rect 282 98 337 100
rect 339 98 340 100
rect 279 97 340 98
rect 144 65 284 69
rect 111 56 236 60
rect 12 51 203 52
rect 12 49 14 51
rect 16 49 103 51
rect 105 49 196 51
rect 198 49 200 51
rect 202 49 203 51
rect 12 48 203 49
rect 232 51 236 56
rect 280 54 284 65
rect 280 52 281 54
rect 283 52 284 54
rect 280 51 284 52
rect 232 49 233 51
rect 235 49 236 51
rect 232 47 236 49
rect 304 50 356 51
rect 304 48 305 50
rect 307 48 356 50
rect 304 47 356 48
rect 352 45 353 47
rect 355 45 356 47
rect 352 44 356 45
rect 159 42 348 43
rect 33 40 74 41
rect 33 38 35 40
rect 37 38 71 40
rect 73 38 74 40
rect 159 40 160 42
rect 162 40 345 42
rect 347 40 348 42
rect 159 39 348 40
rect 367 42 372 105
rect 367 40 368 42
rect 370 40 372 42
rect 33 37 74 38
rect 367 35 372 40
rect 191 34 225 35
rect 191 32 192 34
rect 194 32 222 34
rect 224 32 225 34
rect 191 31 225 32
rect 324 34 372 35
rect 324 32 325 34
rect 327 32 372 34
rect 324 31 372 32
rect 2 16 4 18
rect 6 16 7 18
rect -152 12 -148 15
rect 2 14 7 16
rect -171 8 -148 12
<< alu3 >>
rect 310 117 314 118
rect 310 115 311 117
rect 313 115 314 117
rect -135 99 -131 100
rect -135 97 -134 99
rect -132 97 -131 99
rect -135 76 -131 97
rect 310 76 314 115
rect -250 72 -131 76
rect 195 72 314 76
rect -250 33 -246 72
rect 195 51 199 72
rect 195 49 196 51
rect 198 49 199 51
rect 195 48 199 49
rect -250 31 -249 33
rect -247 31 -246 33
rect -250 30 -246 31
<< alu4 >>
rect 336 98 340 102
rect -276 46 -272 50
<< ptie >>
rect -307 82 -289 84
rect -307 80 -305 82
rect -303 80 -293 82
rect -291 80 -289 82
rect -307 78 -289 80
rect -13 82 -7 84
rect -13 80 -11 82
rect -9 80 -7 82
rect -13 78 -7 80
rect 73 82 99 84
rect 73 80 75 82
rect 77 80 95 82
rect 97 80 99 82
rect 73 78 99 80
rect 296 83 330 85
rect 296 81 298 83
rect 300 81 326 83
rect 328 81 330 83
rect 296 79 330 81
rect 337 83 343 85
rect 337 81 339 83
rect 341 81 343 83
rect 337 79 343 81
rect -279 67 -273 69
rect -279 65 -277 67
rect -275 65 -273 67
rect -279 63 -273 65
rect -266 67 -232 69
rect -266 65 -264 67
rect -262 65 -236 67
rect -234 65 -232 67
rect -266 63 -232 65
rect -35 68 -9 70
rect -35 66 -33 68
rect -31 66 -13 68
rect -11 66 -9 68
rect -35 64 -9 66
rect 71 68 77 70
rect 71 66 73 68
rect 75 66 77 68
rect 71 64 77 66
rect 353 68 371 70
rect 353 66 355 68
rect 357 66 367 68
rect 369 66 371 68
rect 353 64 371 66
<< ntie >>
rect -307 142 -289 144
rect -307 140 -305 142
rect -303 140 -293 142
rect -291 140 -289 142
rect -307 138 -289 140
rect -13 142 -7 144
rect -13 140 -11 142
rect -9 140 -7 142
rect -13 138 -7 140
rect 55 142 61 144
rect 55 140 57 142
rect 59 140 61 142
rect 104 143 110 145
rect 104 141 106 143
rect 108 141 110 143
rect 55 138 61 140
rect 104 139 110 141
rect 220 143 226 145
rect 220 141 222 143
rect 224 141 226 143
rect 220 139 226 141
rect 284 143 290 145
rect 284 141 286 143
rect 288 141 290 143
rect 284 139 290 141
rect 296 143 302 145
rect 296 141 298 143
rect 300 141 302 143
rect 337 143 371 145
rect 296 139 302 141
rect 337 141 339 143
rect 341 141 353 143
rect 355 141 367 143
rect 369 141 371 143
rect 337 139 371 141
rect -307 7 -273 9
rect -307 5 -305 7
rect -303 5 -291 7
rect -289 5 -277 7
rect -275 5 -273 7
rect -238 7 -232 9
rect -307 3 -273 5
rect -238 5 -236 7
rect -234 5 -232 7
rect -238 3 -232 5
rect -226 7 -220 9
rect -226 5 -224 7
rect -222 5 -220 7
rect -226 3 -220 5
rect -162 7 -156 9
rect -162 5 -160 7
rect -158 5 -156 7
rect -162 3 -156 5
rect -46 7 -40 9
rect 3 8 9 10
rect -46 5 -44 7
rect -42 5 -40 7
rect -46 3 -40 5
rect 3 6 5 8
rect 7 6 9 8
rect 3 4 9 6
rect 71 8 77 10
rect 71 6 73 8
rect 75 6 77 8
rect 71 4 77 6
rect 353 8 371 10
rect 353 6 355 8
rect 357 6 367 8
rect 369 6 371 8
rect 353 4 371 6
<< nmos >>
rect -297 92 -295 101
rect -277 87 -275 96
rect -267 87 -265 95
rect -260 87 -258 95
rect -250 87 -248 95
rect -243 87 -241 95
rect -233 89 -231 95
rect -213 81 -211 94
rect -203 84 -201 94
rect -193 87 -191 101
rect -183 87 -181 101
rect -163 81 -161 101
rect -156 81 -154 101
rect -145 81 -143 95
rect -124 81 -122 94
rect -114 84 -112 94
rect -104 87 -102 101
rect -94 87 -92 101
rect -74 81 -72 101
rect -67 81 -65 101
rect -35 95 -33 101
rect -25 95 -23 101
rect -56 81 -54 95
rect -15 92 -13 101
rect 80 94 82 100
rect 90 94 92 100
rect 9 87 11 93
rect 19 87 21 93
rect 26 87 28 93
rect 36 87 38 93
rect 43 87 45 93
rect 53 87 55 93
rect 110 88 112 94
rect 120 88 122 94
rect 127 88 129 94
rect 137 88 139 94
rect 144 88 146 94
rect 154 88 156 94
rect 174 88 176 94
rect 184 88 186 94
rect 191 88 193 94
rect 201 88 203 94
rect 208 88 210 94
rect 218 88 220 94
rect 238 88 240 94
rect 248 88 250 94
rect 255 88 257 94
rect 265 88 267 94
rect 272 88 274 94
rect 282 88 284 94
rect 302 91 304 97
rect 312 91 314 97
rect 322 91 324 97
rect 343 91 345 97
rect 355 85 357 94
rect 362 85 364 94
rect -300 54 -298 63
rect -293 54 -291 63
rect -281 51 -279 57
rect -260 51 -258 57
rect -250 51 -248 57
rect -240 51 -238 57
rect -220 54 -218 60
rect -210 54 -208 60
rect -203 54 -201 60
rect -193 54 -191 60
rect -186 54 -184 60
rect -176 54 -174 60
rect -156 54 -154 60
rect -146 54 -144 60
rect -139 54 -137 60
rect -129 54 -127 60
rect -122 54 -120 60
rect -112 54 -110 60
rect -92 54 -90 60
rect -82 54 -80 60
rect -75 54 -73 60
rect -65 54 -63 60
rect -58 54 -56 60
rect -48 54 -46 60
rect 9 55 11 61
rect 19 55 21 61
rect 26 55 28 61
rect 36 55 38 61
rect 43 55 45 61
rect 53 55 55 61
rect -28 48 -26 54
rect -18 48 -16 54
rect 77 47 79 56
rect 118 53 120 67
rect 87 47 89 53
rect 97 47 99 53
rect 129 47 131 67
rect 136 47 138 67
rect 156 47 158 61
rect 166 47 168 61
rect 176 54 178 64
rect 186 54 188 67
rect 207 53 209 67
rect 218 47 220 67
rect 225 47 227 67
rect 245 47 247 61
rect 255 47 257 61
rect 265 54 267 64
rect 275 54 277 67
rect 295 53 297 59
rect 305 53 307 61
rect 312 53 314 61
rect 322 53 324 61
rect 329 53 331 61
rect 339 52 341 61
rect 359 47 361 56
<< pmos >>
rect -297 113 -295 131
rect -277 123 -275 141
rect -267 125 -265 141
rect -260 125 -258 141
rect -250 125 -248 141
rect -243 125 -241 141
rect -233 113 -231 121
rect -213 116 -211 141
rect -200 116 -198 129
rect -190 113 -188 138
rect -183 113 -181 138
rect -165 113 -163 141
rect -155 113 -153 141
rect -145 113 -143 141
rect -124 116 -122 141
rect -111 116 -109 129
rect -101 113 -99 138
rect -94 113 -92 138
rect -76 113 -74 141
rect -66 113 -64 141
rect -56 113 -54 141
rect -35 120 -33 141
rect -28 120 -26 141
rect -15 113 -13 131
rect 9 121 11 133
rect 19 121 21 133
rect 26 121 28 133
rect 36 121 38 133
rect 43 121 45 133
rect 82 121 84 141
rect 89 121 91 141
rect 53 113 55 119
rect 120 122 122 134
rect 127 122 129 134
rect 137 122 139 134
rect 144 122 146 134
rect 154 122 156 134
rect 174 122 176 134
rect 184 122 186 134
rect 191 122 193 134
rect 201 122 203 134
rect 208 122 210 134
rect 110 114 112 120
rect 238 122 240 134
rect 248 122 250 134
rect 255 122 257 134
rect 265 122 267 134
rect 272 122 274 134
rect 218 114 220 120
rect 302 121 304 133
rect 315 124 317 142
rect 322 124 324 142
rect 282 114 284 120
rect 343 114 345 126
rect 353 114 355 124
rect 363 114 365 124
rect -301 24 -299 34
rect -291 24 -289 34
rect -281 22 -279 34
rect -220 28 -218 34
rect -260 6 -258 24
rect -253 6 -251 24
rect -240 15 -238 27
rect -156 28 -154 34
rect -210 14 -208 26
rect -203 14 -201 26
rect -193 14 -191 26
rect -186 14 -184 26
rect -176 14 -174 26
rect -48 28 -46 34
rect -146 14 -144 26
rect -139 14 -137 26
rect -129 14 -127 26
rect -122 14 -120 26
rect -112 14 -110 26
rect -92 14 -90 26
rect -82 14 -80 26
rect -75 14 -73 26
rect -65 14 -63 26
rect -58 14 -56 26
rect 9 29 11 35
rect -27 7 -25 27
rect -20 7 -18 27
rect 19 15 21 27
rect 26 15 28 27
rect 36 15 38 27
rect 43 15 45 27
rect 53 15 55 27
rect 77 17 79 35
rect 90 7 92 28
rect 97 7 99 28
rect 118 7 120 35
rect 128 7 130 35
rect 138 7 140 35
rect 156 10 158 35
rect 163 10 165 35
rect 173 19 175 32
rect 186 7 188 32
rect 207 7 209 35
rect 217 7 219 35
rect 227 7 229 35
rect 245 10 247 35
rect 252 10 254 35
rect 262 19 264 32
rect 275 7 277 32
rect 295 27 297 35
rect 305 7 307 23
rect 312 7 314 23
rect 322 7 324 23
rect 329 7 331 23
rect 339 7 341 25
rect 359 17 361 35
<< polyct0 >>
rect -251 116 -249 118
rect -276 101 -274 103
rect -258 100 -256 102
rect -205 109 -203 111
rect -211 99 -209 101
rect -155 106 -153 108
rect -145 106 -143 108
rect -116 109 -114 111
rect -122 99 -120 101
rect -66 106 -64 108
rect -56 106 -54 108
rect -17 106 -15 108
rect 35 114 37 116
rect 10 98 12 100
rect 28 98 30 100
rect 128 115 130 117
rect 135 99 137 101
rect 200 115 202 117
rect 153 99 155 101
rect 175 99 177 101
rect 193 99 195 101
rect 264 115 266 117
rect 239 99 241 101
rect 257 99 259 101
rect 304 108 306 110
rect 345 107 347 109
rect -283 39 -281 41
rect -242 38 -240 40
rect -195 47 -193 49
rect -177 47 -175 49
rect -202 31 -200 33
rect -131 47 -129 49
rect -113 47 -111 49
rect -91 47 -89 49
rect -138 31 -136 33
rect -73 47 -71 49
rect -66 31 -64 33
rect 34 48 36 50
rect 52 48 54 50
rect 27 32 29 34
rect 79 40 81 42
rect 118 40 120 42
rect 128 40 130 42
rect 184 47 186 49
rect 178 37 180 39
rect 207 40 209 42
rect 217 40 219 42
rect 273 47 275 49
rect 267 37 269 39
rect 320 46 322 48
rect 338 45 340 47
rect 313 30 315 32
<< polyct1 >>
rect -228 126 -226 128
rect -299 106 -297 108
rect -268 111 -266 113
rect -241 106 -239 108
rect -191 106 -189 108
rect -172 106 -170 108
rect -165 106 -163 108
rect -37 113 -35 115
rect -102 106 -100 108
rect -83 106 -81 108
rect -76 106 -74 108
rect 58 124 60 126
rect -27 106 -25 108
rect 18 108 20 110
rect 105 125 107 127
rect 81 114 83 116
rect 45 106 47 108
rect 223 125 225 127
rect 91 105 93 107
rect 118 107 120 109
rect 145 109 147 111
rect 183 109 185 111
rect 287 125 289 127
rect 210 107 212 109
rect 247 109 249 111
rect 355 131 357 133
rect 274 107 276 109
rect 314 115 316 117
rect 324 107 326 109
rect 364 99 366 101
rect -302 47 -300 49
rect -262 39 -260 41
rect -252 31 -250 33
rect -212 39 -210 41
rect -293 15 -291 17
rect -185 37 -183 39
rect -148 39 -146 41
rect -225 21 -223 23
rect -121 37 -119 39
rect -83 37 -81 39
rect -56 39 -54 41
rect -29 41 -27 43
rect -161 21 -159 23
rect 17 40 19 42
rect -19 32 -17 34
rect -43 21 -41 23
rect 44 38 46 40
rect 89 40 91 42
rect 4 22 6 24
rect 138 40 140 42
rect 145 40 147 42
rect 164 40 166 42
rect 99 33 101 35
rect 227 40 229 42
rect 234 40 236 42
rect 253 40 255 42
rect 303 40 305 42
rect 330 35 332 37
rect 361 40 363 42
rect 290 20 292 22
<< ndifct0 >>
rect -306 94 -304 96
rect -272 89 -270 91
rect -255 89 -253 91
rect -238 91 -236 93
rect -228 91 -226 93
rect -208 86 -206 88
rect -198 89 -196 91
rect -188 97 -186 99
rect -178 97 -176 99
rect -178 90 -176 92
rect -168 90 -166 92
rect -151 83 -149 85
rect -119 86 -117 88
rect -109 89 -107 91
rect -99 97 -97 99
rect -89 97 -87 99
rect -89 90 -87 92
rect -79 90 -77 92
rect -30 97 -28 99
rect -62 83 -60 85
rect 74 96 76 98
rect 95 96 97 98
rect -40 84 -38 86
rect 14 89 16 91
rect 31 89 33 91
rect 48 89 50 91
rect 58 89 60 91
rect 105 90 107 92
rect 115 90 117 92
rect 132 90 134 92
rect 149 90 151 92
rect 179 90 181 92
rect 196 90 198 92
rect 213 90 215 92
rect 223 90 225 92
rect 243 90 245 92
rect 260 90 262 92
rect 277 90 279 92
rect 287 90 289 92
rect 307 93 309 95
rect 317 93 319 95
rect 327 93 329 95
rect -21 84 -19 86
rect 367 90 369 92
rect -305 56 -303 58
rect 83 62 85 64
rect -265 53 -263 55
rect -255 53 -253 55
rect -245 53 -243 55
rect -225 56 -223 58
rect -215 56 -213 58
rect -198 56 -196 58
rect -181 56 -179 58
rect -161 56 -159 58
rect -151 56 -149 58
rect -134 56 -132 58
rect -117 56 -115 58
rect -87 56 -85 58
rect -70 56 -68 58
rect -53 56 -51 58
rect -43 56 -41 58
rect 4 57 6 59
rect 14 57 16 59
rect 31 57 33 59
rect 48 57 50 59
rect 102 62 104 64
rect -33 50 -31 52
rect -12 50 -10 52
rect 124 63 126 65
rect 92 49 94 51
rect 141 56 143 58
rect 151 56 153 58
rect 151 49 153 51
rect 161 49 163 51
rect 171 57 173 59
rect 181 60 183 62
rect 213 63 215 65
rect 230 56 232 58
rect 240 56 242 58
rect 240 49 242 51
rect 250 49 252 51
rect 260 57 262 59
rect 270 60 272 62
rect 290 55 292 57
rect 300 55 302 57
rect 317 57 319 59
rect 334 57 336 59
rect 368 52 370 54
<< ndifct1 >>
rect -292 97 -290 99
rect -282 92 -280 94
rect -218 90 -216 92
rect -140 90 -138 92
rect -129 90 -127 92
rect -51 90 -49 92
rect -10 97 -8 99
rect 85 96 87 98
rect 4 89 6 91
rect 159 90 161 92
rect 169 90 171 92
rect 233 90 235 92
rect 297 93 299 95
rect 338 93 340 95
rect 349 81 351 83
rect -287 65 -285 67
rect -276 53 -274 55
rect -235 53 -233 55
rect -171 56 -169 58
rect -107 56 -105 58
rect -97 56 -95 58
rect 58 57 60 59
rect -23 50 -21 52
rect 72 49 74 51
rect 113 56 115 58
rect 191 56 193 58
rect 202 56 204 58
rect 280 56 282 58
rect 344 54 346 56
rect 354 49 356 51
<< ntiect1 >>
rect -305 140 -303 142
rect -293 140 -291 142
rect -11 140 -9 142
rect 57 140 59 142
rect 106 141 108 143
rect 222 141 224 143
rect 286 141 288 143
rect 298 141 300 143
rect 339 141 341 143
rect 353 141 355 143
rect 367 141 369 143
rect -305 5 -303 7
rect -291 5 -289 7
rect -277 5 -275 7
rect -236 5 -234 7
rect -224 5 -222 7
rect -160 5 -158 7
rect -44 5 -42 7
rect 5 6 7 8
rect 73 6 75 8
rect 355 6 357 8
rect 367 6 369 8
<< ptiect1 >>
rect -305 80 -303 82
rect -293 80 -291 82
rect -11 80 -9 82
rect 75 80 77 82
rect 95 80 97 82
rect 298 81 300 83
rect 326 81 328 83
rect 339 81 341 83
rect -277 65 -275 67
rect -264 65 -262 67
rect -236 65 -234 67
rect -33 66 -31 68
rect -13 66 -11 68
rect 73 66 75 68
rect 355 66 357 68
rect 367 66 369 68
<< pdifct0 >>
rect -303 130 -301 132
rect -272 137 -270 139
rect -255 127 -253 129
rect -238 137 -236 139
rect -228 115 -226 117
rect -207 137 -205 139
rect -195 118 -193 120
rect -172 137 -170 139
rect -172 130 -170 132
rect -160 129 -158 131
rect -160 122 -158 124
rect -150 137 -148 139
rect -150 130 -148 132
rect -118 137 -116 139
rect -106 118 -104 120
rect -83 137 -81 139
rect -83 130 -81 132
rect -71 129 -69 131
rect -71 122 -69 124
rect -61 137 -59 139
rect -61 130 -59 132
rect -40 130 -38 132
rect -21 137 -19 139
rect 14 129 16 131
rect 31 123 33 125
rect 48 129 50 131
rect 96 137 98 139
rect 309 138 311 140
rect 96 130 98 132
rect 115 130 117 132
rect 58 115 60 117
rect 132 124 134 126
rect 149 130 151 132
rect 179 130 181 132
rect 196 124 198 126
rect 213 130 215 132
rect 105 116 107 118
rect 243 130 245 132
rect 260 124 262 126
rect 277 130 279 132
rect 223 116 225 118
rect 327 131 329 133
rect 287 116 289 118
rect 348 116 350 118
rect 358 116 360 118
rect 368 120 370 122
rect -306 26 -304 28
rect -296 30 -294 32
rect -286 30 -284 32
rect -225 30 -223 32
rect -265 15 -263 17
rect -161 30 -159 32
rect -215 16 -213 18
rect -198 22 -196 24
rect -181 16 -179 18
rect -43 30 -41 32
rect -151 16 -149 18
rect -134 22 -132 24
rect -117 16 -115 18
rect -87 16 -85 18
rect -70 22 -68 24
rect 4 31 6 33
rect -53 16 -51 18
rect -34 16 -32 18
rect -247 8 -245 10
rect -34 9 -32 11
rect 14 17 16 19
rect 31 23 33 25
rect 48 17 50 19
rect 83 9 85 11
rect 102 16 104 18
rect 123 16 125 18
rect 123 9 125 11
rect 133 24 135 26
rect 133 17 135 19
rect 145 16 147 18
rect 145 9 147 11
rect 168 28 170 30
rect 180 9 182 11
rect 212 16 214 18
rect 212 9 214 11
rect 222 24 224 26
rect 222 17 224 19
rect 234 16 236 18
rect 234 9 236 11
rect 257 28 259 30
rect 269 9 271 11
rect 290 31 292 33
rect 300 9 302 11
rect 317 19 319 21
rect 334 9 336 11
rect 365 16 367 18
<< pdifct1 >>
rect -282 130 -280 132
rect -292 122 -290 124
rect -292 115 -290 117
rect -218 125 -216 127
rect -218 118 -216 120
rect -140 122 -138 124
rect -140 115 -138 117
rect -129 125 -127 127
rect -129 118 -127 120
rect -51 122 -49 124
rect -51 115 -49 117
rect -10 127 -8 129
rect -10 120 -8 122
rect 4 123 6 125
rect 77 131 79 133
rect 159 124 161 126
rect 169 124 171 126
rect 233 124 235 126
rect 297 129 299 131
rect 338 116 340 118
rect -276 30 -274 32
rect -235 17 -233 19
rect -171 22 -169 24
rect -107 22 -105 24
rect -97 22 -95 24
rect -15 15 -13 17
rect 58 23 60 25
rect 72 26 74 28
rect 72 19 74 21
rect 113 31 115 33
rect 113 24 115 26
rect 191 28 193 30
rect 191 21 193 23
rect 202 31 204 33
rect 202 24 204 26
rect 280 28 282 30
rect 280 21 282 23
rect 354 31 356 33
rect 354 24 356 26
rect 344 16 346 18
<< alu0 >>
rect -305 132 -299 139
rect -274 137 -272 139
rect -270 137 -268 139
rect -274 136 -268 137
rect -239 137 -238 139
rect -236 137 -235 139
rect -239 135 -235 137
rect -209 137 -207 139
rect -205 137 -203 139
rect -209 136 -203 137
rect -174 137 -172 139
rect -170 137 -168 139
rect -305 130 -303 132
rect -301 130 -299 132
rect -305 129 -299 130
rect -264 129 -251 130
rect -293 113 -292 120
rect -307 96 -303 98
rect -307 94 -306 96
rect -304 94 -303 96
rect -293 95 -292 101
rect -307 83 -303 94
rect -264 127 -255 129
rect -253 127 -251 129
rect -264 126 -251 127
rect -276 122 -260 126
rect -276 105 -272 122
rect -174 132 -168 137
rect -152 137 -150 139
rect -148 137 -146 139
rect -174 130 -172 132
rect -170 130 -168 132
rect -174 129 -168 130
rect -161 131 -157 133
rect -161 129 -160 131
rect -158 129 -157 131
rect -152 132 -146 137
rect -120 137 -118 139
rect -116 137 -114 139
rect -120 136 -114 137
rect -85 137 -83 139
rect -81 137 -79 139
rect -152 130 -150 132
rect -148 130 -146 132
rect -152 129 -146 130
rect -85 132 -79 137
rect -63 137 -61 139
rect -59 137 -57 139
rect -85 130 -83 132
rect -81 130 -79 132
rect -85 129 -79 130
rect -72 131 -68 133
rect -72 129 -71 131
rect -69 129 -68 131
rect -63 132 -57 137
rect -23 137 -21 139
rect -19 137 -17 139
rect -23 136 -17 137
rect -63 130 -61 132
rect -59 130 -57 132
rect -63 129 -57 130
rect -42 132 -25 133
rect -42 130 -40 132
rect -38 130 -25 132
rect -42 129 -25 130
rect -204 125 -180 129
rect -161 125 -157 129
rect -252 118 -248 120
rect -269 109 -268 115
rect -252 116 -251 118
rect -249 117 -224 118
rect -249 116 -228 117
rect -252 115 -228 116
rect -226 115 -224 117
rect -252 114 -224 115
rect -277 103 -272 105
rect -252 104 -248 114
rect -277 101 -276 103
rect -274 101 -272 103
rect -259 102 -248 104
rect -277 99 -262 101
rect -276 97 -262 99
rect -259 100 -258 102
rect -256 100 -248 102
rect -259 98 -248 100
rect -273 91 -269 93
rect -273 89 -272 91
rect -270 89 -269 91
rect -273 83 -269 89
rect -266 92 -262 97
rect -228 94 -224 114
rect -240 93 -234 94
rect -266 91 -251 92
rect -266 89 -255 91
rect -253 89 -251 91
rect -266 88 -251 89
rect -240 91 -238 93
rect -236 91 -234 93
rect -240 83 -234 91
rect -230 93 -224 94
rect -230 91 -228 93
rect -226 91 -224 93
rect -230 90 -224 91
rect -206 121 -200 125
rect -184 124 -144 125
rect -184 122 -160 124
rect -158 122 -144 124
rect -206 111 -202 121
rect -196 120 -192 122
rect -184 121 -144 122
rect -196 118 -195 120
rect -193 118 -192 120
rect -196 117 -192 118
rect -206 109 -205 111
rect -203 109 -202 111
rect -206 107 -202 109
rect -199 113 -192 117
rect -199 102 -195 113
rect -156 108 -152 113
rect -156 106 -155 108
rect -153 106 -152 108
rect -213 101 -195 102
rect -213 99 -211 101
rect -209 100 -195 101
rect -209 99 -184 100
rect -213 98 -188 99
rect -199 97 -188 98
rect -186 97 -184 99
rect -199 96 -184 97
rect -179 99 -175 101
rect -179 97 -178 99
rect -176 97 -175 99
rect -179 92 -175 97
rect -156 104 -152 106
rect -148 110 -144 121
rect -148 108 -142 110
rect -148 106 -145 108
rect -143 106 -142 108
rect -148 104 -142 106
rect -148 101 -144 104
rect -164 97 -144 101
rect -164 93 -160 97
rect -200 91 -178 92
rect -209 88 -205 90
rect -200 89 -198 91
rect -196 90 -178 91
rect -176 90 -175 92
rect -196 89 -175 90
rect -170 92 -160 93
rect -170 90 -168 92
rect -166 90 -160 92
rect -170 89 -160 90
rect -115 125 -91 129
rect -72 125 -68 129
rect -117 121 -111 125
rect -95 124 -55 125
rect -95 122 -71 124
rect -69 122 -55 124
rect -117 111 -113 121
rect -107 120 -103 122
rect -95 121 -55 122
rect -107 118 -106 120
rect -104 118 -103 120
rect -107 117 -103 118
rect -117 109 -116 111
rect -114 109 -113 111
rect -117 107 -113 109
rect -110 113 -103 117
rect -110 102 -106 113
rect -67 108 -63 113
rect -67 106 -66 108
rect -64 106 -63 108
rect -124 101 -106 102
rect -124 99 -122 101
rect -120 100 -106 101
rect -120 99 -95 100
rect -124 98 -99 99
rect -110 97 -99 98
rect -97 97 -95 99
rect -110 96 -95 97
rect -90 99 -86 101
rect -90 97 -89 99
rect -87 97 -86 99
rect -90 92 -86 97
rect -67 104 -63 106
rect -59 110 -55 121
rect -29 125 -25 129
rect -29 121 -14 125
rect -59 108 -53 110
rect -59 106 -56 108
rect -54 106 -53 108
rect -59 104 -53 106
rect -59 101 -55 104
rect -75 97 -55 101
rect -75 93 -71 97
rect -39 112 -33 113
rect -18 108 -14 121
rect -11 118 -10 129
rect 12 131 18 139
rect 12 129 14 131
rect 16 129 18 131
rect 12 128 18 129
rect 46 131 52 139
rect 95 137 96 139
rect 98 137 99 139
rect 46 129 48 131
rect 50 129 52 131
rect 46 128 52 129
rect -18 106 -17 108
rect -15 106 -14 108
rect -18 100 -14 106
rect -32 99 -14 100
rect -32 97 -30 99
rect -28 97 -14 99
rect -32 96 -14 97
rect 29 125 35 126
rect 18 123 31 125
rect 33 123 35 125
rect 18 121 35 123
rect 95 132 99 137
rect 95 130 96 132
rect 98 130 99 132
rect -111 91 -89 92
rect -200 88 -175 89
rect -120 88 -116 90
rect -111 89 -109 91
rect -107 90 -89 91
rect -87 90 -86 92
rect -107 89 -86 90
rect -81 92 -71 93
rect -81 90 -79 92
rect -77 90 -71 92
rect -81 89 -71 90
rect 18 118 22 121
rect 9 114 22 118
rect 34 117 62 118
rect 9 100 13 114
rect 34 116 58 117
rect 34 114 35 116
rect 37 115 58 116
rect 60 115 62 117
rect 37 114 62 115
rect 34 102 38 114
rect 27 100 38 102
rect 9 98 10 100
rect 12 98 24 100
rect 9 96 24 98
rect 27 98 28 100
rect 30 98 38 100
rect 27 96 38 98
rect -111 88 -86 89
rect 13 91 17 93
rect 13 89 14 91
rect 16 89 17 91
rect -209 86 -208 88
rect -206 86 -205 88
rect -120 86 -119 88
rect -117 86 -116 88
rect -42 86 -36 87
rect -209 83 -205 86
rect -153 85 -147 86
rect -153 83 -151 85
rect -149 83 -147 85
rect -120 83 -116 86
rect -64 85 -58 86
rect -64 83 -62 85
rect -60 83 -58 85
rect -42 84 -40 86
rect -38 84 -36 86
rect -42 83 -36 84
rect -23 86 -17 87
rect -23 84 -21 86
rect -19 84 -17 86
rect -23 83 -17 84
rect 13 83 17 89
rect 20 92 24 96
rect 58 92 62 114
rect 95 128 99 130
rect 113 132 119 140
rect 113 130 115 132
rect 117 130 119 132
rect 113 129 119 130
rect 147 132 153 140
rect 147 130 149 132
rect 151 130 153 132
rect 147 129 153 130
rect 177 132 183 140
rect 177 130 179 132
rect 181 130 183 132
rect 177 129 183 130
rect 211 132 217 140
rect 211 130 213 132
rect 215 130 217 132
rect 211 129 217 130
rect 241 132 247 140
rect 241 130 243 132
rect 245 130 247 132
rect 241 129 247 130
rect 275 132 281 140
rect 307 138 309 140
rect 311 138 313 140
rect 307 137 313 138
rect 275 130 277 132
rect 279 130 281 132
rect 275 129 281 130
rect 130 126 136 127
rect 130 124 132 126
rect 134 124 147 126
rect 130 122 147 124
rect 143 119 147 122
rect 103 118 131 119
rect 103 116 105 118
rect 107 117 131 118
rect 107 116 128 117
rect 103 115 128 116
rect 130 115 131 117
rect 20 91 35 92
rect 20 89 31 91
rect 33 89 35 91
rect 20 88 35 89
rect 46 91 52 92
rect 46 89 48 91
rect 50 89 52 91
rect 46 83 52 89
rect 56 91 62 92
rect 56 89 58 91
rect 60 89 62 91
rect 56 88 62 89
rect 73 98 77 100
rect 73 96 74 98
rect 76 96 77 98
rect 73 84 77 96
rect 94 98 99 100
rect 94 96 95 98
rect 97 96 99 98
rect 94 94 99 96
rect 95 84 99 94
rect 103 93 107 115
rect 127 103 131 115
rect 143 115 156 119
rect 127 101 138 103
rect 152 101 156 115
rect 127 99 135 101
rect 137 99 138 101
rect 127 97 138 99
rect 141 99 153 101
rect 155 99 156 101
rect 141 97 156 99
rect 141 93 145 97
rect 103 92 109 93
rect 103 90 105 92
rect 107 90 109 92
rect 103 89 109 90
rect 113 92 119 93
rect 113 90 115 92
rect 117 90 119 92
rect 113 84 119 90
rect 130 92 145 93
rect 130 90 132 92
rect 134 90 145 92
rect 130 89 145 90
rect 148 92 152 94
rect 148 90 149 92
rect 151 90 152 92
rect 148 84 152 90
rect 194 126 200 127
rect 183 124 196 126
rect 198 124 200 126
rect 183 122 200 124
rect 258 126 264 127
rect 247 124 260 126
rect 262 124 264 126
rect 247 122 264 124
rect 311 133 331 134
rect 311 131 327 133
rect 329 131 331 133
rect 311 130 331 131
rect 183 119 187 122
rect 174 115 187 119
rect 199 118 227 119
rect 174 101 178 115
rect 199 117 223 118
rect 199 115 200 117
rect 202 116 223 117
rect 225 116 227 118
rect 202 115 227 116
rect 199 103 203 115
rect 192 101 203 103
rect 174 99 175 101
rect 177 99 189 101
rect 174 97 189 99
rect 192 99 193 101
rect 195 99 203 101
rect 192 97 203 99
rect 178 92 182 94
rect 178 90 179 92
rect 181 90 182 92
rect 178 84 182 90
rect 185 93 189 97
rect 223 93 227 115
rect 185 92 200 93
rect 185 90 196 92
rect 198 90 200 92
rect 185 89 200 90
rect 211 92 217 93
rect 211 90 213 92
rect 215 90 217 92
rect 211 84 217 90
rect 221 92 227 93
rect 221 90 223 92
rect 225 90 227 92
rect 221 89 227 90
rect 247 119 251 122
rect 238 115 251 119
rect 263 118 291 119
rect 238 101 242 115
rect 263 117 287 118
rect 263 115 264 117
rect 266 116 287 117
rect 289 116 291 118
rect 266 115 291 116
rect 263 103 267 115
rect 256 101 267 103
rect 238 99 239 101
rect 241 99 253 101
rect 238 97 253 99
rect 256 99 257 101
rect 259 99 267 101
rect 256 97 267 99
rect 242 92 246 94
rect 242 90 243 92
rect 245 90 246 92
rect 242 84 246 90
rect 249 93 253 97
rect 287 93 291 115
rect 249 92 264 93
rect 249 90 260 92
rect 262 90 264 92
rect 249 89 264 90
rect 275 92 281 93
rect 275 90 277 92
rect 279 90 281 92
rect 275 84 281 90
rect 285 92 291 93
rect 285 90 287 92
rect 289 90 291 92
rect 285 89 291 90
rect 299 127 300 130
rect 311 126 315 130
rect 303 122 315 126
rect 303 110 307 122
rect 303 108 304 110
rect 306 108 307 110
rect 303 103 307 108
rect 303 99 320 103
rect 305 95 311 96
rect 305 93 307 95
rect 309 93 311 95
rect 305 84 311 93
rect 316 95 320 99
rect 340 114 341 120
rect 344 119 348 140
rect 367 122 371 140
rect 367 120 368 122
rect 370 120 371 122
rect 344 118 352 119
rect 344 116 348 118
rect 350 116 352 118
rect 344 115 352 116
rect 356 118 362 119
rect 367 118 371 120
rect 356 116 358 118
rect 360 116 362 118
rect 356 110 362 116
rect 343 109 362 110
rect 343 107 345 109
rect 347 107 362 109
rect 343 106 362 107
rect 316 93 317 95
rect 319 93 320 95
rect 316 91 320 93
rect 325 95 331 96
rect 325 93 327 95
rect 329 93 331 95
rect 325 84 331 93
rect 340 95 341 97
rect 352 93 356 106
rect 352 92 371 93
rect 352 90 367 92
rect 369 90 371 92
rect 352 89 371 90
rect -307 58 -288 59
rect -307 56 -305 58
rect -303 56 -288 58
rect -307 55 -288 56
rect -292 42 -288 55
rect -277 51 -276 53
rect -267 55 -261 64
rect -267 53 -265 55
rect -263 53 -261 55
rect -267 52 -261 53
rect -256 55 -252 57
rect -256 53 -255 55
rect -253 53 -252 55
rect -298 41 -279 42
rect -298 39 -283 41
rect -281 39 -279 41
rect -298 38 -279 39
rect -298 32 -292 38
rect -298 30 -296 32
rect -294 30 -292 32
rect -307 28 -303 30
rect -298 29 -292 30
rect -288 32 -280 33
rect -288 30 -286 32
rect -284 30 -280 32
rect -288 29 -280 30
rect -307 26 -306 28
rect -304 26 -303 28
rect -307 8 -303 26
rect -284 8 -280 29
rect -277 28 -276 34
rect -256 49 -252 53
rect -247 55 -241 64
rect -247 53 -245 55
rect -243 53 -241 55
rect -247 52 -241 53
rect -256 45 -239 49
rect -243 40 -239 45
rect -243 38 -242 40
rect -240 38 -239 40
rect -243 26 -239 38
rect -251 22 -239 26
rect -251 18 -247 22
rect -236 18 -235 21
rect -227 58 -221 59
rect -227 56 -225 58
rect -223 56 -221 58
rect -227 55 -221 56
rect -217 58 -211 64
rect -217 56 -215 58
rect -213 56 -211 58
rect -217 55 -211 56
rect -200 58 -185 59
rect -200 56 -198 58
rect -196 56 -185 58
rect -200 55 -185 56
rect -227 33 -223 55
rect -189 51 -185 55
rect -182 58 -178 64
rect -182 56 -181 58
rect -179 56 -178 58
rect -182 54 -178 56
rect -203 49 -192 51
rect -203 47 -195 49
rect -193 47 -192 49
rect -189 49 -174 51
rect -189 47 -177 49
rect -175 47 -174 49
rect -203 45 -192 47
rect -203 33 -199 45
rect -227 32 -202 33
rect -227 30 -225 32
rect -223 31 -202 32
rect -200 31 -199 33
rect -223 30 -199 31
rect -178 33 -174 47
rect -227 29 -199 30
rect -187 29 -174 33
rect -187 26 -183 29
rect -163 58 -157 59
rect -163 56 -161 58
rect -159 56 -157 58
rect -163 55 -157 56
rect -153 58 -147 64
rect -153 56 -151 58
rect -149 56 -147 58
rect -153 55 -147 56
rect -136 58 -121 59
rect -136 56 -134 58
rect -132 56 -121 58
rect -136 55 -121 56
rect -163 33 -159 55
rect -125 51 -121 55
rect -118 58 -114 64
rect -118 56 -117 58
rect -115 56 -114 58
rect -118 54 -114 56
rect -139 49 -128 51
rect -139 47 -131 49
rect -129 47 -128 49
rect -125 49 -110 51
rect -125 47 -113 49
rect -111 47 -110 49
rect -139 45 -128 47
rect -139 33 -135 45
rect -163 32 -138 33
rect -163 30 -161 32
rect -159 31 -138 32
rect -136 31 -135 33
rect -159 30 -135 31
rect -114 33 -110 47
rect -163 29 -135 30
rect -123 29 -110 33
rect -123 26 -119 29
rect -267 17 -247 18
rect -267 15 -265 17
rect -263 15 -247 17
rect -267 14 -247 15
rect -200 24 -183 26
rect -200 22 -198 24
rect -196 22 -183 24
rect -200 21 -194 22
rect -136 24 -119 26
rect -136 22 -134 24
rect -132 22 -119 24
rect -136 21 -130 22
rect -88 58 -84 64
rect -88 56 -87 58
rect -85 56 -84 58
rect -88 54 -84 56
rect -81 58 -66 59
rect -81 56 -70 58
rect -68 56 -66 58
rect -81 55 -66 56
rect -55 58 -49 64
rect -55 56 -53 58
rect -51 56 -49 58
rect -55 55 -49 56
rect -45 58 -39 59
rect -45 56 -43 58
rect -41 56 -39 58
rect -45 55 -39 56
rect -81 51 -77 55
rect -92 49 -77 51
rect -92 47 -91 49
rect -89 47 -77 49
rect -74 49 -63 51
rect -74 47 -73 49
rect -71 47 -63 49
rect -92 33 -88 47
rect -74 45 -63 47
rect -92 29 -79 33
rect -67 33 -63 45
rect -43 33 -39 55
rect -35 54 -31 64
rect -35 52 -30 54
rect -35 50 -33 52
rect -31 50 -30 52
rect -35 48 -30 50
rect -13 52 -9 64
rect -13 50 -12 52
rect -10 50 -9 52
rect -13 48 -9 50
rect 2 59 8 60
rect 2 57 4 59
rect 6 57 8 59
rect 2 56 8 57
rect 12 59 18 65
rect 12 57 14 59
rect 16 57 18 59
rect 12 56 18 57
rect 29 59 44 60
rect 29 57 31 59
rect 33 57 44 59
rect 29 56 44 57
rect -67 31 -66 33
rect -64 32 -39 33
rect -64 31 -43 32
rect -67 30 -43 31
rect -41 30 -39 32
rect -67 29 -39 30
rect -83 26 -79 29
rect -83 24 -66 26
rect -83 22 -70 24
rect -68 22 -66 24
rect -72 21 -66 22
rect -217 18 -211 19
rect -217 16 -215 18
rect -213 16 -211 18
rect -249 10 -243 11
rect -249 8 -247 10
rect -245 8 -243 10
rect -217 8 -211 16
rect -183 18 -177 19
rect -183 16 -181 18
rect -179 16 -177 18
rect -183 8 -177 16
rect -153 18 -147 19
rect -153 16 -151 18
rect -149 16 -147 18
rect -153 8 -147 16
rect -119 18 -113 19
rect -119 16 -117 18
rect -115 16 -113 18
rect -119 8 -113 16
rect -89 18 -83 19
rect -89 16 -87 18
rect -85 16 -83 18
rect -89 8 -83 16
rect -55 18 -49 19
rect -55 16 -53 18
rect -51 16 -49 18
rect -55 8 -49 16
rect -35 18 -31 20
rect 2 34 6 56
rect 40 52 44 56
rect 47 59 51 65
rect 81 64 87 65
rect 81 62 83 64
rect 85 62 87 64
rect 81 61 87 62
rect 100 64 106 65
rect 100 62 102 64
rect 104 62 106 64
rect 122 63 124 65
rect 126 63 128 65
rect 122 62 128 63
rect 180 62 184 65
rect 211 63 213 65
rect 215 63 217 65
rect 211 62 217 63
rect 269 62 273 65
rect 100 61 106 62
rect 180 60 181 62
rect 183 60 184 62
rect 269 60 270 62
rect 272 60 273 62
rect 47 57 48 59
rect 50 57 51 59
rect 47 55 51 57
rect 150 59 175 60
rect 26 50 37 52
rect 26 48 34 50
rect 36 48 37 50
rect 40 50 55 52
rect 40 48 52 50
rect 54 48 55 50
rect 26 46 37 48
rect 26 34 30 46
rect 2 33 27 34
rect 2 31 4 33
rect 6 32 27 33
rect 29 32 30 34
rect 6 31 30 32
rect 51 34 55 48
rect 2 30 30 31
rect 42 30 55 34
rect 42 27 46 30
rect 135 58 145 59
rect 135 56 141 58
rect 143 56 145 58
rect 135 55 145 56
rect 150 58 171 59
rect 150 56 151 58
rect 153 57 171 58
rect 173 57 175 59
rect 180 58 184 60
rect 239 59 264 60
rect 153 56 175 57
rect -35 16 -34 18
rect -32 16 -31 18
rect -35 11 -31 16
rect 29 25 46 27
rect 29 23 31 25
rect 33 23 46 25
rect 29 22 35 23
rect 78 51 96 52
rect 78 49 92 51
rect 94 49 96 51
rect 78 48 96 49
rect 78 42 82 48
rect 78 40 79 42
rect 81 40 82 42
rect 12 19 18 20
rect 12 17 14 19
rect 16 17 18 19
rect -35 9 -34 11
rect -32 9 -31 11
rect 12 9 18 17
rect 46 19 52 20
rect 46 17 48 19
rect 50 17 52 19
rect 46 9 52 17
rect 74 19 75 30
rect 78 27 82 40
rect 97 35 103 36
rect 135 51 139 55
rect 119 47 139 51
rect 119 44 123 47
rect 117 42 123 44
rect 117 40 118 42
rect 120 40 123 42
rect 117 38 123 40
rect 78 23 93 27
rect 89 19 93 23
rect 119 27 123 38
rect 127 42 131 44
rect 150 51 154 56
rect 150 49 151 51
rect 153 49 154 51
rect 150 47 154 49
rect 159 51 174 52
rect 159 49 161 51
rect 163 50 174 51
rect 163 49 188 50
rect 159 48 184 49
rect 170 47 184 48
rect 186 47 188 49
rect 170 46 188 47
rect 127 40 128 42
rect 130 40 131 42
rect 127 35 131 40
rect 170 35 174 46
rect 167 31 174 35
rect 177 39 181 41
rect 177 37 178 39
rect 180 37 181 39
rect 167 30 171 31
rect 167 28 168 30
rect 170 28 171 30
rect 119 26 159 27
rect 167 26 171 28
rect 177 27 181 37
rect 119 24 133 26
rect 135 24 159 26
rect 119 23 159 24
rect 175 23 181 27
rect 132 19 136 23
rect 155 19 179 23
rect 224 58 234 59
rect 224 56 230 58
rect 232 56 234 58
rect 224 55 234 56
rect 239 58 260 59
rect 239 56 240 58
rect 242 57 260 58
rect 262 57 264 59
rect 269 58 273 60
rect 242 56 264 57
rect 224 51 228 55
rect 208 47 228 51
rect 208 44 212 47
rect 206 42 212 44
rect 206 40 207 42
rect 209 40 212 42
rect 206 38 212 40
rect 208 27 212 38
rect 216 42 220 44
rect 239 51 243 56
rect 239 49 240 51
rect 242 49 243 51
rect 239 47 243 49
rect 248 51 263 52
rect 248 49 250 51
rect 252 50 263 51
rect 252 49 277 50
rect 248 48 273 49
rect 259 47 273 48
rect 275 47 277 49
rect 259 46 277 47
rect 216 40 217 42
rect 219 40 220 42
rect 216 35 220 40
rect 259 35 263 46
rect 256 31 263 35
rect 266 39 270 41
rect 266 37 267 39
rect 269 37 270 39
rect 256 30 260 31
rect 256 28 257 30
rect 259 28 260 30
rect 208 26 248 27
rect 256 26 260 28
rect 266 27 270 37
rect 208 24 222 26
rect 224 24 248 26
rect 208 23 248 24
rect 264 23 270 27
rect 288 57 294 58
rect 288 55 290 57
rect 292 55 294 57
rect 288 54 294 55
rect 298 57 304 65
rect 298 55 300 57
rect 302 55 304 57
rect 315 59 330 60
rect 315 57 317 59
rect 319 57 330 59
rect 315 56 330 57
rect 298 54 304 55
rect 288 34 292 54
rect 326 51 330 56
rect 333 59 337 65
rect 333 57 334 59
rect 336 57 337 59
rect 333 55 337 57
rect 312 48 323 50
rect 312 46 320 48
rect 322 46 323 48
rect 326 49 340 51
rect 326 47 341 49
rect 312 44 323 46
rect 336 45 338 47
rect 340 45 341 47
rect 312 34 316 44
rect 336 43 341 45
rect 288 33 316 34
rect 288 31 290 33
rect 292 32 316 33
rect 292 31 313 32
rect 288 30 313 31
rect 315 30 316 32
rect 332 33 333 39
rect 312 28 316 30
rect 221 19 225 23
rect 244 19 268 23
rect 89 18 106 19
rect 89 16 102 18
rect 104 16 106 18
rect 89 15 106 16
rect 121 18 127 19
rect 121 16 123 18
rect 125 16 127 18
rect 81 11 87 12
rect 81 9 83 11
rect 85 9 87 11
rect 121 11 127 16
rect 132 17 133 19
rect 135 17 136 19
rect 132 15 136 17
rect 143 18 149 19
rect 143 16 145 18
rect 147 16 149 18
rect 121 9 123 11
rect 125 9 127 11
rect 143 11 149 16
rect 210 18 216 19
rect 210 16 212 18
rect 214 16 216 18
rect 143 9 145 11
rect 147 9 149 11
rect 178 11 184 12
rect 178 9 180 11
rect 182 9 184 11
rect 210 11 216 16
rect 221 17 222 19
rect 224 17 225 19
rect 221 15 225 17
rect 232 18 238 19
rect 232 16 234 18
rect 236 16 238 18
rect 210 9 212 11
rect 214 9 216 11
rect 232 11 238 16
rect 336 26 340 43
rect 324 22 340 26
rect 315 21 328 22
rect 315 19 317 21
rect 319 19 328 21
rect 367 54 371 65
rect 356 47 357 53
rect 367 52 368 54
rect 370 52 371 54
rect 367 50 371 52
rect 356 28 357 35
rect 315 18 328 19
rect 363 18 369 19
rect 363 16 365 18
rect 367 16 369 18
rect 232 9 234 11
rect 236 9 238 11
rect 267 11 273 12
rect 267 9 269 11
rect 271 9 273 11
rect 299 11 303 13
rect 299 9 300 11
rect 302 9 303 11
rect 332 11 338 12
rect 332 9 334 11
rect 336 9 338 11
rect 363 9 369 16
<< via1 >>
rect -306 106 -304 108
rect -291 101 -289 103
rect -283 106 -281 108
rect -263 114 -261 116
rect -243 98 -241 100
rect -160 114 -158 116
rect -219 94 -217 96
rect -171 97 -169 99
rect -138 97 -136 99
rect -130 114 -128 116
rect -98 106 -96 108
rect 58 130 60 132
rect -9 108 -7 110
rect -41 97 -39 99
rect 27 108 29 110
rect 48 97 50 99
rect 104 130 106 132
rect 224 129 226 131
rect 288 130 290 132
rect 89 123 91 125
rect 73 111 75 113
rect 97 115 99 117
rect 117 99 119 101
rect 140 108 142 110
rect 160 108 162 110
rect 188 108 190 110
rect 212 99 214 101
rect 232 99 234 101
rect 257 111 259 113
rect 280 98 282 100
rect 296 111 298 113
rect 320 124 322 126
rect 328 107 330 109
rect 353 124 355 126
rect 369 107 371 109
rect 337 98 339 100
rect -275 48 -273 50
rect -307 39 -305 41
rect -291 22 -289 24
rect -266 39 -264 41
rect -258 22 -256 24
rect -234 35 -232 37
rect -218 48 -216 50
rect -195 35 -193 37
rect -170 47 -168 49
rect -150 47 -148 49
rect -126 38 -124 40
rect -98 38 -96 40
rect -78 38 -76 40
rect -55 47 -53 49
rect -35 31 -33 33
rect -11 35 -9 37
rect -27 23 -25 25
rect -226 16 -224 18
rect -162 17 -160 19
rect -42 16 -40 18
rect 14 49 16 51
rect 35 38 37 40
rect 103 49 105 51
rect 71 38 73 40
rect 4 16 6 18
rect 160 40 162 42
rect 192 32 194 34
rect 200 49 202 51
rect 233 49 235 51
rect 281 52 283 54
rect 222 32 224 34
rect 305 48 307 50
rect 325 32 327 34
rect 345 40 347 42
rect 353 45 355 47
rect 368 40 370 42
<< via2 >>
rect -134 97 -132 99
rect 311 115 313 117
rect -249 31 -247 33
rect 196 49 198 51
<< labels >>
rlabel alu1 198 69 198 69 5 Vss
rlabel alu1 346 27 346 27 5 b_test
rlabel alu1 301 49 301 49 5 Bn
rlabel alu1 290 15 290 15 5 Binv
rlabel alu1 282 38 282 38 5 Sum
rlabel via1 326 33 326 33 5 B
rlabel alu1 145 51 145 51 5 A
rlabel alu1 198 5 198 5 5 Vdd
rlabel alu1 234 49 234 49 5 Cin
rlabel alu1 60 37 60 37 1 COUT
rlabel alu1 32 5 32 5 2 vdd
rlabel alu1 32 69 32 69 2 vss
rlabel alu1 72 36 72 36 1 fafs_cout
rlabel via1 15 50 15 50 1 in1
rlabel alu2 40 38 40 38 1 in2
rlabel alu1 145 108 145 108 4 a0
rlabel alu1 133 80 133 80 4 vss
rlabel alu1 121 104 121 104 4 a1
rlabel alu1 133 144 133 144 4 vdd
rlabel via1 161 108 161 108 1 y0
rlabel alu1 197 80 197 80 6 vss
rlabel alu1 197 144 197 144 6 vdd
rlabel alu2 210 100 210 100 1 k1
rlabel alu1 232 107 233 109 1 y1
rlabel alu1 277 100 277 100 1 a3
rlabel alu1 261 144 261 144 6 vdd
rlabel alu1 261 80 261 80 6 vss
rlabel alu1 113 100 113 100 4 a1
rlabel alu1 354 128 354 128 6 a
rlabel alu1 362 100 362 100 6 b
rlabel alu1 362 132 362 132 6 a
rlabel alu1 354 144 354 144 6 vdd
rlabel alu1 169 105 169 105 1 out
rlabel alu1 313 80 313 80 6 vss
rlabel alu1 313 116 313 116 6 a
rlabel alu1 313 144 313 144 6 vdd
rlabel alu1 321 108 321 108 6 b
rlabel alu1 321 124 321 124 6 a
rlabel space 293 79 333 147 1 or
rlabel space 335 79 375 147 1 and
rlabel alu1 329 112 329 112 6 b
rlabel alu4 338 99 338 99 1 z3
rlabel via1 297 112 297 112 1 z2
rlabel space 96 79 293 147 1 4x1_mux
rlabel via1 188 110 188 110 1 k0
rlabel alu1 370 104 370 104 6 b
rlabel alu1 354 80 354 80 6 vss
rlabel space 65 1 376 77 1 fafs
rlabel space 0 1 64 77 1 shift_mux
rlabel alu1 4 17 4 17 3 fafs_en
rlabel alu1 74 119 74 119 6 z
rlabel alu1 82 99 82 99 6 z
rlabel alu1 86 79 86 79 6 vss
rlabel alu1 86 143 86 143 6 vdd
rlabel alu1 94 107 94 107 1 l1
rlabel alu1 85 119 85 119 1 l0
rlabel ab 71 78 100 147 1 decoder
rlabel alu1 252 109 252 109 1 or_out
rlabel alu1 224 134 224 134 1 s1
rlabel alu2 163 131 163 131 1 s0
rlabel alu1 -134 79 -134 79 1 Vss
rlabel alu1 -282 121 -282 121 1 b_test
rlabel alu1 -237 99 -237 99 1 Bn
rlabel alu1 -226 133 -226 133 1 Binv
rlabel alu1 -218 110 -218 110 1 Sum
rlabel via1 -262 115 -262 115 1 B
rlabel alu1 -81 97 -81 97 1 A
rlabel alu1 -134 143 -134 143 1 Vdd
rlabel alu1 -170 99 -170 99 1 Cin
rlabel alu1 4 111 4 111 5 COUT
rlabel alu1 32 143 32 143 6 vdd
rlabel alu1 32 79 32 79 6 vss
rlabel alu1 -8 112 -8 112 5 fafs_cout
rlabel via1 49 98 49 98 5 in1
rlabel alu2 24 110 24 110 5 in2
rlabel alu1 -81 40 -81 40 8 a0
rlabel alu1 -69 68 -69 68 8 vss
rlabel alu1 -57 44 -57 44 8 a1
rlabel alu1 -69 4 -69 4 8 vdd
rlabel via1 -97 40 -97 40 5 y0
rlabel alu1 -133 68 -133 68 2 vss
rlabel alu1 -133 4 -133 4 2 vdd
rlabel alu2 -146 48 -146 48 5 k1
rlabel alu1 -169 39 -168 41 5 y1
rlabel alu1 -213 48 -213 48 5 a3
rlabel alu1 -197 4 -197 4 2 vdd
rlabel alu1 -197 68 -197 68 2 vss
rlabel alu1 -49 48 -49 48 8 a1
rlabel alu1 -290 20 -290 20 2 a
rlabel alu1 -298 48 -298 48 2 b
rlabel alu1 -298 16 -298 16 2 a
rlabel alu1 -290 4 -290 4 2 vdd
rlabel alu1 -105 43 -105 43 5 out
rlabel alu1 -249 68 -249 68 2 vss
rlabel alu1 -249 32 -249 32 2 a
rlabel alu1 -249 4 -249 4 2 vdd
rlabel alu1 -257 40 -257 40 2 b
rlabel alu1 -257 24 -257 24 2 a
rlabel space -269 1 -229 69 5 or
rlabel space -311 1 -271 69 5 and
rlabel alu1 -265 36 -265 36 2 b
rlabel alu4 -274 49 -274 49 5 z3
rlabel via1 -233 36 -233 36 5 z2
rlabel space -229 1 -32 69 5 4x1_mux
rlabel via1 -124 38 -124 38 5 k0
rlabel alu1 -306 44 -306 44 2 b
rlabel alu1 -290 68 -290 68 2 vss
rlabel space -312 71 -1 147 5 fafs
rlabel space 0 71 64 147 5 shift_mux
rlabel alu1 60 131 60 131 7 fafs_en
rlabel alu1 -10 29 -10 29 2 z
rlabel alu1 -18 49 -18 49 2 z
rlabel alu1 -22 69 -22 69 2 vss
rlabel alu1 -22 5 -22 5 2 vdd
rlabel alu1 -30 41 -30 41 5 l1
rlabel alu1 -21 29 -21 29 5 l0
rlabel ab -36 1 -7 70 5 decoder
rlabel alu1 -188 39 -188 39 5 or_out
rlabel alu1 -160 14 -160 14 5 s1
rlabel alu2 -99 17 -99 17 5 s0
<< end >>
