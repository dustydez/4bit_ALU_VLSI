magic
tech scmos
timestamp 1760387970
<< ab >>
rect 157 74 266 146
rect 268 74 310 146
rect 312 74 375 146
rect 382 76 412 146
rect 413 145 490 146
rect 497 145 603 146
rect 609 145 686 146
rect 413 77 645 145
rect 646 77 686 145
rect 377 74 409 76
rect 279 70 311 72
rect 2 1 42 69
rect 43 1 275 69
rect 2 0 79 1
rect 85 0 191 1
rect 198 0 275 1
rect 276 0 306 70
rect 313 0 376 72
rect 378 0 420 72
rect 422 0 531 72
<< nwell >>
rect 0 107 688 146
rect 0 106 382 107
rect 308 39 336 40
rect 375 39 688 40
rect 0 0 688 39
<< pwell >>
rect 382 106 688 107
rect 0 66 688 106
rect 0 40 316 66
rect 336 40 688 66
rect 0 39 308 40
rect 336 39 375 40
<< poly >>
rect 35 140 37 144
rect 45 140 47 144
rect 52 140 54 144
rect 62 140 64 144
rect 69 140 71 144
rect 99 140 101 144
rect 15 130 17 135
rect 82 127 88 129
rect 82 125 84 127
rect 86 125 88 127
rect 15 109 17 112
rect 11 107 17 109
rect 11 105 13 107
rect 15 105 17 107
rect 11 103 17 105
rect 35 104 37 122
rect 45 114 47 124
rect 42 112 48 114
rect 42 110 44 112
rect 46 110 48 112
rect 42 108 48 110
rect 52 109 54 124
rect 62 119 64 124
rect 59 117 65 119
rect 59 115 61 117
rect 63 115 65 117
rect 59 113 65 115
rect 69 109 71 124
rect 79 123 88 125
rect 79 120 81 123
rect 122 137 124 142
rect 129 137 131 142
rect 147 140 149 144
rect 157 140 159 144
rect 167 140 169 144
rect 188 140 190 144
rect 112 128 114 133
rect 15 100 17 103
rect 34 102 40 104
rect 34 100 36 102
rect 38 100 40 102
rect 34 98 40 100
rect 35 95 37 98
rect 15 86 17 91
rect 45 94 47 108
rect 52 107 64 109
rect 52 101 58 103
rect 52 99 54 101
rect 56 99 58 101
rect 52 97 58 99
rect 52 94 54 97
rect 62 94 64 107
rect 69 107 75 109
rect 69 105 71 107
rect 73 105 75 107
rect 69 103 75 105
rect 69 94 71 103
rect 79 94 81 112
rect 99 102 101 115
rect 112 112 114 115
rect 211 137 213 142
rect 218 137 220 142
rect 236 140 238 144
rect 246 140 248 144
rect 256 140 258 144
rect 277 140 279 144
rect 284 140 286 144
rect 201 128 203 133
rect 105 110 114 112
rect 105 108 107 110
rect 109 108 111 110
rect 122 109 124 112
rect 129 109 131 112
rect 147 109 149 112
rect 157 109 159 112
rect 167 109 169 112
rect 105 106 111 108
rect 99 100 105 102
rect 99 98 101 100
rect 103 98 105 100
rect 99 96 105 98
rect 99 93 101 96
rect 109 93 111 106
rect 119 107 125 109
rect 119 105 121 107
rect 123 105 125 107
rect 119 103 125 105
rect 129 107 151 109
rect 129 105 140 107
rect 142 105 147 107
rect 149 105 151 107
rect 129 103 151 105
rect 155 107 161 109
rect 155 105 157 107
rect 159 105 161 107
rect 155 103 161 105
rect 165 107 171 109
rect 165 105 167 107
rect 169 105 171 107
rect 165 103 171 105
rect 119 100 121 103
rect 129 100 131 103
rect 149 100 151 103
rect 156 100 158 103
rect 35 81 37 86
rect 45 81 47 86
rect 52 81 54 86
rect 62 78 64 86
rect 69 82 71 86
rect 79 78 81 88
rect 62 76 81 78
rect 99 76 101 80
rect 109 78 111 83
rect 119 81 121 86
rect 129 81 131 86
rect 167 94 169 103
rect 188 102 190 115
rect 201 112 203 115
rect 394 140 396 144
rect 401 140 403 144
rect 297 130 299 135
rect 321 132 323 137
rect 331 132 333 137
rect 338 132 340 137
rect 348 132 350 137
rect 355 132 357 137
rect 277 116 279 119
rect 273 114 279 116
rect 273 112 275 114
rect 277 112 279 114
rect 194 110 203 112
rect 194 108 196 110
rect 198 108 200 110
rect 211 109 213 112
rect 218 109 220 112
rect 236 109 238 112
rect 246 109 248 112
rect 256 109 258 112
rect 273 110 279 112
rect 194 106 200 108
rect 188 100 194 102
rect 188 98 190 100
rect 192 98 194 100
rect 188 96 194 98
rect 188 93 190 96
rect 198 93 200 106
rect 208 107 214 109
rect 208 105 210 107
rect 212 105 214 107
rect 208 103 214 105
rect 218 107 240 109
rect 218 105 229 107
rect 231 105 236 107
rect 238 105 240 107
rect 218 103 240 105
rect 244 107 250 109
rect 244 105 246 107
rect 248 105 250 107
rect 244 103 250 105
rect 254 107 260 109
rect 254 105 256 107
rect 258 105 260 107
rect 254 103 260 105
rect 208 100 210 103
rect 218 100 220 103
rect 238 100 240 103
rect 245 100 247 103
rect 149 76 151 80
rect 156 76 158 80
rect 167 76 169 80
rect 188 76 190 80
rect 198 78 200 83
rect 208 81 210 86
rect 218 81 220 86
rect 256 94 258 103
rect 277 100 279 110
rect 284 109 286 119
rect 368 125 374 127
rect 368 123 370 125
rect 372 123 374 125
rect 297 109 299 112
rect 283 107 289 109
rect 283 105 285 107
rect 287 105 289 107
rect 283 103 289 105
rect 293 107 299 109
rect 293 105 295 107
rect 297 105 299 107
rect 293 103 299 105
rect 287 100 289 103
rect 297 100 299 103
rect 321 101 323 120
rect 331 111 333 120
rect 328 109 334 111
rect 328 107 330 109
rect 332 107 334 109
rect 328 105 334 107
rect 338 107 340 120
rect 348 117 350 120
rect 345 115 351 117
rect 345 113 347 115
rect 349 113 351 115
rect 345 111 351 113
rect 355 109 357 120
rect 365 121 374 123
rect 365 118 367 121
rect 627 141 629 145
rect 634 141 636 145
rect 432 133 434 138
rect 439 133 441 138
rect 449 133 451 138
rect 456 133 458 138
rect 466 133 468 138
rect 486 133 488 138
rect 496 133 498 138
rect 503 133 505 138
rect 513 133 515 138
rect 520 133 522 138
rect 550 133 552 138
rect 560 133 562 138
rect 567 133 569 138
rect 577 133 579 138
rect 584 133 586 138
rect 415 126 421 128
rect 415 124 417 126
rect 419 124 421 126
rect 415 122 424 124
rect 394 117 396 120
rect 391 115 397 117
rect 391 113 393 115
rect 395 113 397 115
rect 355 107 361 109
rect 338 105 350 107
rect 277 89 279 94
rect 287 89 289 94
rect 320 99 326 101
rect 320 97 322 99
rect 324 97 326 99
rect 320 95 326 97
rect 321 92 323 95
rect 331 92 333 105
rect 338 99 344 101
rect 338 97 340 99
rect 342 97 344 99
rect 338 95 344 97
rect 338 92 340 95
rect 348 92 350 105
rect 355 105 357 107
rect 359 105 361 107
rect 355 103 361 105
rect 355 92 357 103
rect 365 92 367 112
rect 391 111 397 113
rect 392 99 394 111
rect 401 108 403 120
rect 422 119 424 122
rect 533 126 539 128
rect 533 124 535 126
rect 537 124 539 126
rect 401 106 407 108
rect 401 104 403 106
rect 405 104 407 106
rect 401 102 407 104
rect 402 99 404 102
rect 422 93 424 113
rect 432 110 434 121
rect 439 118 441 121
rect 438 116 444 118
rect 438 114 440 116
rect 442 114 444 116
rect 438 112 444 114
rect 428 108 434 110
rect 449 108 451 121
rect 456 112 458 121
rect 428 106 430 108
rect 432 106 434 108
rect 428 104 434 106
rect 432 93 434 104
rect 439 106 451 108
rect 455 110 461 112
rect 455 108 457 110
rect 459 108 461 110
rect 455 106 461 108
rect 439 93 441 106
rect 445 100 451 102
rect 445 98 447 100
rect 449 98 451 100
rect 445 96 451 98
rect 449 93 451 96
rect 456 93 458 106
rect 466 102 468 121
rect 486 102 488 121
rect 496 112 498 121
rect 493 110 499 112
rect 493 108 495 110
rect 497 108 499 110
rect 493 106 499 108
rect 503 108 505 121
rect 513 118 515 121
rect 510 116 516 118
rect 510 114 512 116
rect 514 114 516 116
rect 510 112 516 114
rect 520 110 522 121
rect 530 122 539 124
rect 530 119 532 122
rect 614 132 616 136
rect 597 126 603 128
rect 597 124 599 126
rect 601 124 603 126
rect 520 108 526 110
rect 503 106 515 108
rect 463 100 469 102
rect 463 98 465 100
rect 467 98 469 100
rect 463 96 469 98
rect 485 100 491 102
rect 485 98 487 100
rect 489 98 491 100
rect 485 96 491 98
rect 466 93 468 96
rect 486 93 488 96
rect 496 93 498 106
rect 503 100 509 102
rect 503 98 505 100
rect 507 98 509 100
rect 503 96 509 98
rect 503 93 505 96
rect 513 93 515 106
rect 520 106 522 108
rect 524 106 526 108
rect 520 104 526 106
rect 520 93 522 104
rect 530 93 532 113
rect 550 102 552 121
rect 560 112 562 121
rect 557 110 563 112
rect 557 108 559 110
rect 561 108 563 110
rect 557 106 563 108
rect 567 108 569 121
rect 577 118 579 121
rect 574 116 580 118
rect 574 114 576 116
rect 578 114 580 116
rect 574 112 580 114
rect 584 110 586 121
rect 594 122 603 124
rect 594 119 596 122
rect 665 132 671 134
rect 665 130 667 132
rect 669 130 671 132
rect 655 125 657 130
rect 665 128 671 130
rect 584 108 590 110
rect 567 106 579 108
rect 549 100 555 102
rect 549 98 551 100
rect 553 98 555 100
rect 549 96 555 98
rect 550 93 552 96
rect 560 93 562 106
rect 567 100 573 102
rect 567 98 569 100
rect 571 98 573 100
rect 567 96 573 98
rect 567 93 569 96
rect 577 93 579 106
rect 584 106 586 108
rect 588 106 590 108
rect 584 104 590 106
rect 584 93 586 104
rect 594 93 596 113
rect 614 111 616 120
rect 627 118 629 123
rect 624 116 630 118
rect 624 114 626 116
rect 628 114 630 116
rect 624 112 630 114
rect 614 109 620 111
rect 614 107 616 109
rect 618 107 620 109
rect 614 105 620 107
rect 614 96 616 105
rect 624 96 626 112
rect 634 110 636 123
rect 665 123 667 128
rect 675 123 677 128
rect 655 110 657 113
rect 665 110 667 113
rect 634 108 640 110
rect 634 106 636 108
rect 638 106 640 108
rect 634 104 640 106
rect 655 108 661 110
rect 655 106 657 108
rect 659 106 661 108
rect 665 107 669 110
rect 655 104 661 106
rect 634 96 636 104
rect 655 96 657 104
rect 297 86 299 91
rect 392 88 394 93
rect 402 88 404 93
rect 667 93 669 107
rect 675 102 677 113
rect 674 100 680 102
rect 674 98 676 100
rect 678 98 680 100
rect 674 96 680 98
rect 674 93 676 96
rect 321 81 323 86
rect 331 81 333 86
rect 338 81 340 86
rect 238 76 240 80
rect 245 76 247 80
rect 256 76 258 80
rect 348 78 350 86
rect 355 82 357 86
rect 365 78 367 86
rect 348 76 367 78
rect 422 79 424 87
rect 432 83 434 87
rect 439 79 441 87
rect 449 82 451 87
rect 456 82 458 87
rect 466 82 468 87
rect 486 82 488 87
rect 496 82 498 87
rect 503 82 505 87
rect 422 77 441 79
rect 513 79 515 87
rect 520 83 522 87
rect 530 79 532 87
rect 550 82 552 87
rect 560 82 562 87
rect 567 82 569 87
rect 513 77 532 79
rect 577 79 579 87
rect 584 83 586 87
rect 594 79 596 87
rect 614 86 616 90
rect 624 86 626 90
rect 634 86 636 90
rect 655 86 657 90
rect 577 77 596 79
rect 667 79 669 84
rect 674 79 676 84
rect 12 62 14 67
rect 19 62 21 67
rect 92 67 111 69
rect 31 56 33 60
rect 52 56 54 60
rect 62 56 64 60
rect 72 56 74 60
rect 92 59 94 67
rect 102 59 104 63
rect 109 59 111 67
rect 156 67 175 69
rect 119 59 121 64
rect 126 59 128 64
rect 136 59 138 64
rect 156 59 158 67
rect 166 59 168 63
rect 173 59 175 67
rect 247 67 266 69
rect 183 59 185 64
rect 190 59 192 64
rect 200 59 202 64
rect 220 59 222 64
rect 230 59 232 64
rect 237 59 239 64
rect 247 59 249 67
rect 254 59 256 63
rect 264 59 266 67
rect 321 68 340 70
rect 321 60 323 68
rect 331 60 333 64
rect 338 60 340 68
rect 430 66 432 70
rect 441 66 443 70
rect 448 66 450 70
rect 348 60 350 65
rect 355 60 357 65
rect 365 60 367 65
rect 12 50 14 53
rect 8 48 14 50
rect 8 46 10 48
rect 12 46 14 48
rect 8 44 14 46
rect 11 33 13 44
rect 19 39 21 53
rect 284 53 286 58
rect 294 53 296 58
rect 389 55 391 60
rect 31 42 33 50
rect 52 42 54 50
rect 27 40 33 42
rect 19 36 23 39
rect 27 38 29 40
rect 31 38 33 40
rect 27 36 33 38
rect 48 40 54 42
rect 48 38 50 40
rect 52 38 54 40
rect 48 36 54 38
rect 21 33 23 36
rect 31 33 33 36
rect 11 18 13 23
rect 21 18 23 23
rect 52 23 54 36
rect 62 34 64 50
rect 72 41 74 50
rect 68 39 74 41
rect 68 37 70 39
rect 72 37 74 39
rect 68 35 74 37
rect 58 32 64 34
rect 58 30 60 32
rect 62 30 64 32
rect 58 28 64 30
rect 59 23 61 28
rect 72 26 74 35
rect 92 33 94 53
rect 102 42 104 53
rect 98 40 104 42
rect 98 38 100 40
rect 102 38 104 40
rect 109 40 111 53
rect 119 50 121 53
rect 115 48 121 50
rect 115 46 117 48
rect 119 46 121 48
rect 115 44 121 46
rect 126 40 128 53
rect 136 50 138 53
rect 133 48 139 50
rect 133 46 135 48
rect 137 46 139 48
rect 133 44 139 46
rect 109 38 121 40
rect 98 36 104 38
rect 17 16 23 18
rect 31 16 33 21
rect 17 14 19 16
rect 21 14 23 16
rect 17 12 23 14
rect 92 24 94 27
rect 85 22 94 24
rect 102 25 104 36
rect 108 32 114 34
rect 108 30 110 32
rect 112 30 114 32
rect 108 28 114 30
rect 109 25 111 28
rect 119 25 121 38
rect 125 38 131 40
rect 125 36 127 38
rect 129 36 131 38
rect 125 34 131 36
rect 126 25 128 34
rect 136 25 138 44
rect 156 33 158 53
rect 166 42 168 53
rect 162 40 168 42
rect 162 38 164 40
rect 166 38 168 40
rect 173 40 175 53
rect 183 50 185 53
rect 179 48 185 50
rect 179 46 181 48
rect 183 46 185 48
rect 179 44 185 46
rect 190 40 192 53
rect 200 50 202 53
rect 220 50 222 53
rect 197 48 203 50
rect 197 46 199 48
rect 201 46 203 48
rect 197 44 203 46
rect 219 48 225 50
rect 219 46 221 48
rect 223 46 225 48
rect 219 44 225 46
rect 173 38 185 40
rect 162 36 168 38
rect 85 20 87 22
rect 89 20 91 22
rect 85 18 91 20
rect 72 10 74 14
rect 156 24 158 27
rect 149 22 158 24
rect 166 25 168 36
rect 172 32 178 34
rect 172 30 174 32
rect 176 30 178 32
rect 172 28 178 30
rect 173 25 175 28
rect 183 25 185 38
rect 189 38 195 40
rect 189 36 191 38
rect 193 36 195 38
rect 189 34 195 36
rect 190 25 192 34
rect 200 25 202 44
rect 220 25 222 44
rect 230 40 232 53
rect 237 50 239 53
rect 237 48 243 50
rect 237 46 239 48
rect 241 46 243 48
rect 237 44 243 46
rect 247 40 249 53
rect 227 38 233 40
rect 227 36 229 38
rect 231 36 233 38
rect 227 34 233 36
rect 237 38 249 40
rect 254 42 256 53
rect 254 40 260 42
rect 254 38 256 40
rect 258 38 260 40
rect 230 25 232 34
rect 237 25 239 38
rect 254 36 260 38
rect 244 32 250 34
rect 244 30 246 32
rect 248 30 250 32
rect 244 28 250 30
rect 247 25 249 28
rect 254 25 256 36
rect 264 33 266 53
rect 284 44 286 47
rect 281 42 287 44
rect 281 40 283 42
rect 285 40 287 42
rect 281 38 287 40
rect 149 20 151 22
rect 153 20 155 22
rect 149 18 155 20
rect 264 24 266 27
rect 285 26 287 38
rect 294 35 296 47
rect 291 33 297 35
rect 321 34 323 54
rect 331 43 333 54
rect 327 41 333 43
rect 327 39 329 41
rect 331 39 333 41
rect 338 41 340 54
rect 348 51 350 54
rect 344 49 350 51
rect 344 47 346 49
rect 348 47 350 49
rect 344 45 350 47
rect 355 41 357 54
rect 365 51 367 54
rect 362 49 368 51
rect 362 47 364 49
rect 366 47 368 49
rect 362 45 368 47
rect 399 52 401 57
rect 409 52 411 57
rect 338 39 350 41
rect 327 37 333 39
rect 291 31 293 33
rect 295 31 297 33
rect 291 29 297 31
rect 292 26 294 29
rect 264 22 273 24
rect 267 20 269 22
rect 271 20 273 22
rect 267 18 273 20
rect 102 8 104 13
rect 109 8 111 13
rect 119 8 121 13
rect 126 8 128 13
rect 136 8 138 13
rect 166 8 168 13
rect 173 8 175 13
rect 183 8 185 13
rect 190 8 192 13
rect 200 8 202 13
rect 220 8 222 13
rect 230 8 232 13
rect 237 8 239 13
rect 247 8 249 13
rect 254 8 256 13
rect 52 1 54 5
rect 59 1 61 5
rect 321 25 323 28
rect 314 23 323 25
rect 331 26 333 37
rect 337 33 343 35
rect 337 31 339 33
rect 341 31 343 33
rect 337 29 343 31
rect 338 26 340 29
rect 348 26 350 39
rect 354 39 360 41
rect 354 37 356 39
rect 358 37 360 39
rect 354 35 360 37
rect 355 26 357 35
rect 365 26 367 45
rect 389 43 391 46
rect 399 43 401 46
rect 389 41 395 43
rect 389 39 391 41
rect 393 39 395 41
rect 389 37 395 39
rect 399 41 405 43
rect 399 39 401 41
rect 403 39 405 41
rect 399 37 405 39
rect 389 34 391 37
rect 314 21 316 23
rect 318 21 320 23
rect 314 19 320 21
rect 402 27 404 37
rect 409 36 411 46
rect 430 43 432 52
rect 468 60 470 65
rect 478 60 480 65
rect 488 63 490 68
rect 498 66 500 70
rect 519 66 521 70
rect 530 66 532 70
rect 537 66 539 70
rect 441 43 443 46
rect 448 43 450 46
rect 468 43 470 46
rect 478 43 480 46
rect 428 41 434 43
rect 428 39 430 41
rect 432 39 434 41
rect 428 37 434 39
rect 438 41 444 43
rect 438 39 440 41
rect 442 39 444 41
rect 438 37 444 39
rect 448 41 470 43
rect 448 39 450 41
rect 452 39 457 41
rect 459 39 470 41
rect 448 37 470 39
rect 474 41 480 43
rect 474 39 476 41
rect 478 39 480 41
rect 474 37 480 39
rect 488 40 490 53
rect 498 50 500 53
rect 494 48 500 50
rect 494 46 496 48
rect 498 46 500 48
rect 494 44 500 46
rect 488 38 494 40
rect 409 34 415 36
rect 430 34 432 37
rect 440 34 442 37
rect 450 34 452 37
rect 468 34 470 37
rect 475 34 477 37
rect 488 36 490 38
rect 492 36 494 38
rect 485 34 494 36
rect 409 32 411 34
rect 413 32 415 34
rect 409 30 415 32
rect 409 27 411 30
rect 331 9 333 14
rect 338 9 340 14
rect 348 9 350 14
rect 355 9 357 14
rect 365 9 367 14
rect 389 11 391 16
rect 285 2 287 6
rect 292 2 294 6
rect 485 31 487 34
rect 498 31 500 44
rect 519 43 521 52
rect 557 60 559 65
rect 567 60 569 65
rect 577 63 579 68
rect 587 66 589 70
rect 607 68 626 70
rect 607 58 609 68
rect 617 60 619 64
rect 624 60 626 68
rect 634 60 636 65
rect 641 60 643 65
rect 651 60 653 65
rect 530 43 532 46
rect 537 43 539 46
rect 557 43 559 46
rect 567 43 569 46
rect 517 41 523 43
rect 517 39 519 41
rect 521 39 523 41
rect 517 37 523 39
rect 527 41 533 43
rect 527 39 529 41
rect 531 39 533 41
rect 527 37 533 39
rect 537 41 559 43
rect 537 39 539 41
rect 541 39 546 41
rect 548 39 559 41
rect 537 37 559 39
rect 563 41 569 43
rect 563 39 565 41
rect 567 39 569 41
rect 563 37 569 39
rect 577 40 579 53
rect 587 50 589 53
rect 583 48 589 50
rect 583 46 585 48
rect 587 46 589 48
rect 583 44 589 46
rect 577 38 583 40
rect 519 34 521 37
rect 529 34 531 37
rect 539 34 541 37
rect 557 34 559 37
rect 564 34 566 37
rect 577 36 579 38
rect 581 36 583 38
rect 574 34 583 36
rect 485 13 487 18
rect 402 2 404 6
rect 409 2 411 6
rect 430 2 432 6
rect 440 2 442 6
rect 450 2 452 6
rect 468 4 470 9
rect 475 4 477 9
rect 574 31 576 34
rect 587 31 589 44
rect 607 34 609 52
rect 617 43 619 52
rect 613 41 619 43
rect 613 39 615 41
rect 617 39 619 41
rect 613 37 619 39
rect 624 39 626 52
rect 634 49 636 52
rect 630 47 636 49
rect 630 45 632 47
rect 634 45 636 47
rect 630 43 636 45
rect 624 37 636 39
rect 641 38 643 52
rect 671 55 673 60
rect 651 48 653 51
rect 648 46 654 48
rect 648 44 650 46
rect 652 44 654 46
rect 648 42 654 44
rect 671 43 673 46
rect 574 13 576 18
rect 498 2 500 6
rect 519 2 521 6
rect 529 2 531 6
rect 539 2 541 6
rect 557 4 559 9
rect 564 4 566 9
rect 607 23 609 26
rect 600 21 609 23
rect 617 22 619 37
rect 623 31 629 33
rect 623 29 625 31
rect 627 29 629 31
rect 623 27 629 29
rect 624 22 626 27
rect 634 22 636 37
rect 640 36 646 38
rect 640 34 642 36
rect 644 34 646 36
rect 640 32 646 34
rect 641 22 643 32
rect 651 24 653 42
rect 671 41 677 43
rect 671 39 673 41
rect 675 39 677 41
rect 671 37 677 39
rect 671 34 673 37
rect 600 19 602 21
rect 604 19 606 21
rect 600 17 606 19
rect 671 11 673 16
rect 587 2 589 6
rect 617 2 619 6
rect 624 2 626 6
rect 634 2 636 6
rect 641 2 643 6
rect 651 2 653 6
<< ndif >>
rect 4 95 15 100
rect 4 93 6 95
rect 8 93 15 95
rect 4 91 15 93
rect 17 98 24 100
rect 17 96 20 98
rect 22 96 24 98
rect 17 94 24 96
rect 17 91 22 94
rect 28 93 35 95
rect 28 91 30 93
rect 32 91 35 93
rect 28 89 35 91
rect 30 86 35 89
rect 37 94 42 95
rect 37 90 45 94
rect 37 88 40 90
rect 42 88 45 90
rect 37 86 45 88
rect 47 86 52 94
rect 54 90 62 94
rect 54 88 57 90
rect 59 88 62 90
rect 54 86 62 88
rect 64 86 69 94
rect 71 92 79 94
rect 71 90 74 92
rect 76 90 79 92
rect 71 88 79 90
rect 81 92 88 94
rect 114 93 119 100
rect 81 90 84 92
rect 86 90 88 92
rect 81 88 88 90
rect 92 91 99 93
rect 92 89 94 91
rect 96 89 99 91
rect 71 86 77 88
rect 92 87 99 89
rect 94 80 99 87
rect 101 87 109 93
rect 101 85 104 87
rect 106 85 109 87
rect 101 83 109 85
rect 111 90 119 93
rect 111 88 114 90
rect 116 88 119 90
rect 111 86 119 88
rect 121 98 129 100
rect 121 96 124 98
rect 126 96 129 98
rect 121 86 129 96
rect 131 98 138 100
rect 131 96 134 98
rect 136 96 138 98
rect 131 91 138 96
rect 144 93 149 100
rect 131 89 134 91
rect 136 89 138 91
rect 131 86 138 89
rect 142 91 149 93
rect 142 89 144 91
rect 146 89 149 91
rect 142 87 149 89
rect 111 83 116 86
rect 101 80 106 83
rect 144 80 149 87
rect 151 80 156 100
rect 158 94 165 100
rect 158 84 167 94
rect 158 82 161 84
rect 163 82 167 84
rect 158 80 167 82
rect 169 91 176 94
rect 203 93 208 100
rect 169 89 172 91
rect 174 89 176 91
rect 169 87 176 89
rect 181 91 188 93
rect 181 89 183 91
rect 185 89 188 91
rect 181 87 188 89
rect 169 80 174 87
rect 183 80 188 87
rect 190 87 198 93
rect 190 85 193 87
rect 195 85 198 87
rect 190 83 198 85
rect 200 90 208 93
rect 200 88 203 90
rect 205 88 208 90
rect 200 86 208 88
rect 210 98 218 100
rect 210 96 213 98
rect 215 96 218 98
rect 210 86 218 96
rect 220 98 227 100
rect 220 96 223 98
rect 225 96 227 98
rect 220 91 227 96
rect 233 93 238 100
rect 220 89 223 91
rect 225 89 227 91
rect 220 86 227 89
rect 231 91 238 93
rect 231 89 233 91
rect 235 89 238 91
rect 231 87 238 89
rect 200 83 205 86
rect 190 80 195 83
rect 233 80 238 87
rect 240 80 245 100
rect 247 94 254 100
rect 270 94 277 100
rect 279 98 287 100
rect 279 96 282 98
rect 284 96 287 98
rect 279 94 287 96
rect 289 94 297 100
rect 247 84 256 94
rect 247 82 250 84
rect 252 82 256 84
rect 247 80 256 82
rect 258 91 265 94
rect 258 89 261 91
rect 263 89 265 91
rect 258 87 265 89
rect 270 87 275 94
rect 291 91 297 94
rect 299 98 306 100
rect 299 96 302 98
rect 304 96 306 98
rect 299 94 306 96
rect 299 91 304 94
rect 384 97 392 99
rect 384 95 386 97
rect 388 95 392 97
rect 384 93 392 95
rect 394 97 402 99
rect 394 95 397 97
rect 399 95 402 97
rect 394 93 402 95
rect 404 97 411 99
rect 404 95 407 97
rect 409 95 411 97
rect 404 93 411 95
rect 607 94 614 96
rect 291 87 295 91
rect 258 80 263 87
rect 270 85 276 87
rect 270 83 272 85
rect 274 83 276 85
rect 270 81 276 83
rect 289 85 295 87
rect 314 90 321 92
rect 314 88 316 90
rect 318 88 321 90
rect 314 86 321 88
rect 323 90 331 92
rect 323 88 326 90
rect 328 88 331 90
rect 323 86 331 88
rect 333 86 338 92
rect 340 90 348 92
rect 340 88 343 90
rect 345 88 348 90
rect 340 86 348 88
rect 350 86 355 92
rect 357 90 365 92
rect 357 88 360 90
rect 362 88 365 90
rect 357 86 365 88
rect 367 90 374 92
rect 367 88 370 90
rect 372 88 374 90
rect 415 91 422 93
rect 415 89 417 91
rect 419 89 422 91
rect 367 86 374 88
rect 415 87 422 89
rect 424 91 432 93
rect 424 89 427 91
rect 429 89 432 91
rect 424 87 432 89
rect 434 87 439 93
rect 441 91 449 93
rect 441 89 444 91
rect 446 89 449 91
rect 441 87 449 89
rect 451 87 456 93
rect 458 91 466 93
rect 458 89 461 91
rect 463 89 466 91
rect 458 87 466 89
rect 468 91 475 93
rect 468 89 471 91
rect 473 89 475 91
rect 468 87 475 89
rect 479 91 486 93
rect 479 89 481 91
rect 483 89 486 91
rect 479 87 486 89
rect 488 91 496 93
rect 488 89 491 91
rect 493 89 496 91
rect 488 87 496 89
rect 498 87 503 93
rect 505 91 513 93
rect 505 89 508 91
rect 510 89 513 91
rect 505 87 513 89
rect 515 87 520 93
rect 522 91 530 93
rect 522 89 525 91
rect 527 89 530 91
rect 522 87 530 89
rect 532 91 539 93
rect 532 89 535 91
rect 537 89 539 91
rect 532 87 539 89
rect 543 91 550 93
rect 543 89 545 91
rect 547 89 550 91
rect 543 87 550 89
rect 552 91 560 93
rect 552 89 555 91
rect 557 89 560 91
rect 552 87 560 89
rect 562 87 567 93
rect 569 91 577 93
rect 569 89 572 91
rect 574 89 577 91
rect 569 87 577 89
rect 579 87 584 93
rect 586 91 594 93
rect 586 89 589 91
rect 591 89 594 91
rect 586 87 594 89
rect 596 91 603 93
rect 596 89 599 91
rect 601 89 603 91
rect 607 92 609 94
rect 611 92 614 94
rect 607 90 614 92
rect 616 94 624 96
rect 616 92 619 94
rect 621 92 624 94
rect 616 90 624 92
rect 626 94 634 96
rect 626 92 629 94
rect 631 92 634 94
rect 626 90 634 92
rect 636 94 643 96
rect 636 92 639 94
rect 641 92 643 94
rect 636 90 643 92
rect 648 94 655 96
rect 648 92 650 94
rect 652 92 655 94
rect 648 90 655 92
rect 657 93 665 96
rect 657 90 667 93
rect 596 87 603 89
rect 289 83 291 85
rect 293 83 295 85
rect 289 81 295 83
rect 659 84 667 90
rect 669 84 674 93
rect 676 91 683 93
rect 676 89 679 91
rect 681 89 683 91
rect 676 87 683 89
rect 676 84 681 87
rect 659 82 665 84
rect 659 80 661 82
rect 663 80 665 82
rect 659 78 665 80
rect 23 66 29 68
rect 23 64 25 66
rect 27 64 29 66
rect 23 62 29 64
rect 7 59 12 62
rect 5 57 12 59
rect 5 55 7 57
rect 9 55 12 57
rect 5 53 12 55
rect 14 53 19 62
rect 21 56 29 62
rect 393 63 399 65
rect 393 61 395 63
rect 397 61 399 63
rect 85 57 92 59
rect 21 53 31 56
rect 23 50 31 53
rect 33 54 40 56
rect 33 52 36 54
rect 38 52 40 54
rect 33 50 40 52
rect 45 54 52 56
rect 45 52 47 54
rect 49 52 52 54
rect 45 50 52 52
rect 54 54 62 56
rect 54 52 57 54
rect 59 52 62 54
rect 54 50 62 52
rect 64 54 72 56
rect 64 52 67 54
rect 69 52 72 54
rect 64 50 72 52
rect 74 54 81 56
rect 74 52 77 54
rect 79 52 81 54
rect 85 55 87 57
rect 89 55 92 57
rect 85 53 92 55
rect 94 57 102 59
rect 94 55 97 57
rect 99 55 102 57
rect 94 53 102 55
rect 104 53 109 59
rect 111 57 119 59
rect 111 55 114 57
rect 116 55 119 57
rect 111 53 119 55
rect 121 53 126 59
rect 128 57 136 59
rect 128 55 131 57
rect 133 55 136 57
rect 128 53 136 55
rect 138 57 145 59
rect 138 55 141 57
rect 143 55 145 57
rect 138 53 145 55
rect 149 57 156 59
rect 149 55 151 57
rect 153 55 156 57
rect 149 53 156 55
rect 158 57 166 59
rect 158 55 161 57
rect 163 55 166 57
rect 158 53 166 55
rect 168 53 173 59
rect 175 57 183 59
rect 175 55 178 57
rect 180 55 183 57
rect 175 53 183 55
rect 185 53 190 59
rect 192 57 200 59
rect 192 55 195 57
rect 197 55 200 57
rect 192 53 200 55
rect 202 57 209 59
rect 202 55 205 57
rect 207 55 209 57
rect 202 53 209 55
rect 213 57 220 59
rect 213 55 215 57
rect 217 55 220 57
rect 213 53 220 55
rect 222 57 230 59
rect 222 55 225 57
rect 227 55 230 57
rect 222 53 230 55
rect 232 53 237 59
rect 239 57 247 59
rect 239 55 242 57
rect 244 55 247 57
rect 239 53 247 55
rect 249 53 254 59
rect 256 57 264 59
rect 256 55 259 57
rect 261 55 264 57
rect 256 53 264 55
rect 266 57 273 59
rect 314 58 321 60
rect 266 55 269 57
rect 271 55 273 57
rect 266 53 273 55
rect 314 56 316 58
rect 318 56 321 58
rect 314 54 321 56
rect 323 58 331 60
rect 323 56 326 58
rect 328 56 331 58
rect 323 54 331 56
rect 333 54 338 60
rect 340 58 348 60
rect 340 56 343 58
rect 345 56 348 58
rect 340 54 348 56
rect 350 54 355 60
rect 357 58 365 60
rect 357 56 360 58
rect 362 56 365 58
rect 357 54 365 56
rect 367 58 374 60
rect 367 56 370 58
rect 372 56 374 58
rect 367 54 374 56
rect 393 59 399 61
rect 412 63 418 65
rect 412 61 414 63
rect 416 61 418 63
rect 412 59 418 61
rect 425 59 430 66
rect 393 55 397 59
rect 74 50 81 52
rect 277 51 284 53
rect 277 49 279 51
rect 281 49 284 51
rect 277 47 284 49
rect 286 51 294 53
rect 286 49 289 51
rect 291 49 294 51
rect 286 47 294 49
rect 296 51 304 53
rect 296 49 300 51
rect 302 49 304 51
rect 296 47 304 49
rect 384 52 389 55
rect 382 50 389 52
rect 382 48 384 50
rect 386 48 389 50
rect 382 46 389 48
rect 391 52 397 55
rect 413 52 418 59
rect 423 57 430 59
rect 423 55 425 57
rect 427 55 430 57
rect 423 52 430 55
rect 432 64 441 66
rect 432 62 436 64
rect 438 62 441 64
rect 432 52 441 62
rect 391 46 399 52
rect 401 50 409 52
rect 401 48 404 50
rect 406 48 409 50
rect 401 46 409 48
rect 411 46 418 52
rect 434 46 441 52
rect 443 46 448 66
rect 450 59 455 66
rect 493 63 498 66
rect 483 60 488 63
rect 450 57 457 59
rect 450 55 453 57
rect 455 55 457 57
rect 450 53 457 55
rect 461 57 468 60
rect 461 55 463 57
rect 465 55 468 57
rect 450 46 455 53
rect 461 50 468 55
rect 461 48 463 50
rect 465 48 468 50
rect 461 46 468 48
rect 470 50 478 60
rect 470 48 473 50
rect 475 48 478 50
rect 470 46 478 48
rect 480 58 488 60
rect 480 56 483 58
rect 485 56 488 58
rect 480 53 488 56
rect 490 61 498 63
rect 490 59 493 61
rect 495 59 498 61
rect 490 53 498 59
rect 500 59 505 66
rect 514 59 519 66
rect 500 57 507 59
rect 500 55 503 57
rect 505 55 507 57
rect 500 53 507 55
rect 512 57 519 59
rect 512 55 514 57
rect 516 55 519 57
rect 480 46 485 53
rect 512 52 519 55
rect 521 64 530 66
rect 521 62 525 64
rect 527 62 530 64
rect 521 52 530 62
rect 523 46 530 52
rect 532 46 537 66
rect 539 59 544 66
rect 582 63 587 66
rect 572 60 577 63
rect 539 57 546 59
rect 539 55 542 57
rect 544 55 546 57
rect 539 53 546 55
rect 550 57 557 60
rect 550 55 552 57
rect 554 55 557 57
rect 539 46 544 53
rect 550 50 557 55
rect 550 48 552 50
rect 554 48 557 50
rect 550 46 557 48
rect 559 50 567 60
rect 559 48 562 50
rect 564 48 567 50
rect 559 46 567 48
rect 569 58 577 60
rect 569 56 572 58
rect 574 56 577 58
rect 569 53 577 56
rect 579 61 587 63
rect 579 59 582 61
rect 584 59 587 61
rect 579 53 587 59
rect 589 59 594 66
rect 589 57 596 59
rect 611 58 617 60
rect 589 55 592 57
rect 594 55 596 57
rect 589 53 596 55
rect 600 56 607 58
rect 600 54 602 56
rect 604 54 607 56
rect 569 46 574 53
rect 600 52 607 54
rect 609 56 617 58
rect 609 54 612 56
rect 614 54 617 56
rect 609 52 617 54
rect 619 52 624 60
rect 626 58 634 60
rect 626 56 629 58
rect 631 56 634 58
rect 626 52 634 56
rect 636 52 641 60
rect 643 58 651 60
rect 643 56 646 58
rect 648 56 651 58
rect 643 52 651 56
rect 646 51 651 52
rect 653 57 658 60
rect 653 55 660 57
rect 653 53 656 55
rect 658 53 660 55
rect 653 51 660 53
rect 666 52 671 55
rect 664 50 671 52
rect 664 48 666 50
rect 668 48 671 50
rect 664 46 671 48
rect 673 53 684 55
rect 673 51 680 53
rect 682 51 684 53
rect 673 46 684 51
<< pdif >>
rect 6 131 13 133
rect 6 129 9 131
rect 11 130 13 131
rect 30 133 35 140
rect 28 131 35 133
rect 11 129 15 130
rect 6 112 15 129
rect 17 125 22 130
rect 28 129 30 131
rect 32 129 35 131
rect 28 127 35 129
rect 17 123 24 125
rect 17 121 20 123
rect 22 121 24 123
rect 30 122 35 127
rect 37 138 45 140
rect 37 136 40 138
rect 42 136 45 138
rect 37 124 45 136
rect 47 124 52 140
rect 54 128 62 140
rect 54 126 57 128
rect 59 126 62 128
rect 54 124 62 126
rect 64 124 69 140
rect 71 138 78 140
rect 71 136 74 138
rect 76 136 78 138
rect 71 128 78 136
rect 71 124 77 128
rect 94 128 99 140
rect 37 122 42 124
rect 17 116 24 121
rect 17 114 20 116
rect 22 114 24 116
rect 17 112 24 114
rect 73 120 77 124
rect 92 126 99 128
rect 92 124 94 126
rect 96 124 99 126
rect 73 112 79 120
rect 81 118 86 120
rect 92 119 99 124
rect 81 116 88 118
rect 81 114 84 116
rect 86 114 88 116
rect 92 117 94 119
rect 96 117 99 119
rect 92 115 99 117
rect 101 138 110 140
rect 101 136 105 138
rect 107 136 110 138
rect 133 138 147 140
rect 133 137 140 138
rect 101 128 110 136
rect 117 128 122 137
rect 101 115 112 128
rect 114 119 122 128
rect 114 117 117 119
rect 119 117 122 119
rect 114 115 122 117
rect 81 112 88 114
rect 117 112 122 115
rect 124 112 129 137
rect 131 136 140 137
rect 142 136 147 138
rect 131 131 147 136
rect 131 129 140 131
rect 142 129 147 131
rect 131 112 147 129
rect 149 130 157 140
rect 149 128 152 130
rect 154 128 157 130
rect 149 123 157 128
rect 149 121 152 123
rect 154 121 157 123
rect 149 112 157 121
rect 159 138 167 140
rect 159 136 162 138
rect 164 136 167 138
rect 159 131 167 136
rect 159 129 162 131
rect 164 129 167 131
rect 159 112 167 129
rect 169 125 174 140
rect 183 128 188 140
rect 181 126 188 128
rect 169 123 176 125
rect 169 121 172 123
rect 174 121 176 123
rect 169 116 176 121
rect 169 114 172 116
rect 174 114 176 116
rect 181 124 183 126
rect 185 124 188 126
rect 181 119 188 124
rect 181 117 183 119
rect 185 117 188 119
rect 181 115 188 117
rect 190 138 199 140
rect 190 136 194 138
rect 196 136 199 138
rect 222 138 236 140
rect 222 137 229 138
rect 190 128 199 136
rect 206 128 211 137
rect 190 115 201 128
rect 203 119 211 128
rect 203 117 206 119
rect 208 117 211 119
rect 203 115 211 117
rect 169 112 176 114
rect 206 112 211 115
rect 213 112 218 137
rect 220 136 229 137
rect 231 136 236 138
rect 220 131 236 136
rect 220 129 229 131
rect 231 129 236 131
rect 220 112 236 129
rect 238 130 246 140
rect 238 128 241 130
rect 243 128 246 130
rect 238 123 246 128
rect 238 121 241 123
rect 243 121 246 123
rect 238 112 246 121
rect 248 138 256 140
rect 248 136 251 138
rect 253 136 256 138
rect 248 131 256 136
rect 248 129 251 131
rect 253 129 256 131
rect 248 112 256 129
rect 258 125 263 140
rect 272 133 277 140
rect 270 131 277 133
rect 270 129 272 131
rect 274 129 277 131
rect 270 127 277 129
rect 258 123 265 125
rect 258 121 261 123
rect 263 121 265 123
rect 258 116 265 121
rect 272 119 277 127
rect 279 119 284 140
rect 286 138 295 140
rect 286 136 291 138
rect 293 136 295 138
rect 286 130 295 136
rect 389 134 394 140
rect 387 132 394 134
rect 286 119 297 130
rect 258 114 261 116
rect 263 114 265 116
rect 258 112 265 114
rect 289 112 297 119
rect 299 128 306 130
rect 299 126 302 128
rect 304 126 306 128
rect 316 126 321 132
rect 299 121 306 126
rect 299 119 302 121
rect 304 119 306 121
rect 314 124 321 126
rect 314 122 316 124
rect 318 122 321 124
rect 314 120 321 122
rect 323 130 331 132
rect 323 128 326 130
rect 328 128 331 130
rect 323 120 331 128
rect 333 120 338 132
rect 340 124 348 132
rect 340 122 343 124
rect 345 122 348 124
rect 340 120 348 122
rect 350 120 355 132
rect 357 130 364 132
rect 357 128 360 130
rect 362 128 364 130
rect 387 130 389 132
rect 391 130 394 132
rect 387 128 394 130
rect 357 126 364 128
rect 357 120 363 126
rect 299 117 306 119
rect 299 112 304 117
rect 359 118 363 120
rect 389 120 394 128
rect 396 120 401 140
rect 403 138 412 140
rect 618 139 627 141
rect 403 136 408 138
rect 410 136 412 138
rect 403 131 412 136
rect 618 137 621 139
rect 623 137 627 139
rect 403 129 408 131
rect 410 129 412 131
rect 403 126 412 129
rect 425 131 432 133
rect 425 129 427 131
rect 429 129 432 131
rect 425 127 432 129
rect 403 120 411 126
rect 359 112 365 118
rect 367 116 374 118
rect 367 114 370 116
rect 372 114 374 116
rect 367 112 374 114
rect 426 121 432 127
rect 434 121 439 133
rect 441 125 449 133
rect 441 123 444 125
rect 446 123 449 125
rect 441 121 449 123
rect 451 121 456 133
rect 458 131 466 133
rect 458 129 461 131
rect 463 129 466 131
rect 458 121 466 129
rect 468 127 473 133
rect 481 127 486 133
rect 468 125 475 127
rect 468 123 471 125
rect 473 123 475 125
rect 468 121 475 123
rect 479 125 486 127
rect 479 123 481 125
rect 483 123 486 125
rect 479 121 486 123
rect 488 131 496 133
rect 488 129 491 131
rect 493 129 496 131
rect 488 121 496 129
rect 498 121 503 133
rect 505 125 513 133
rect 505 123 508 125
rect 510 123 513 125
rect 505 121 513 123
rect 515 121 520 133
rect 522 131 529 133
rect 522 129 525 131
rect 527 129 529 131
rect 522 127 529 129
rect 522 121 528 127
rect 545 127 550 133
rect 426 119 430 121
rect 415 117 422 119
rect 415 115 417 117
rect 419 115 422 117
rect 415 113 422 115
rect 424 113 430 119
rect 524 119 528 121
rect 543 125 550 127
rect 543 123 545 125
rect 547 123 550 125
rect 543 121 550 123
rect 552 131 560 133
rect 552 129 555 131
rect 557 129 560 131
rect 552 121 560 129
rect 562 121 567 133
rect 569 125 577 133
rect 569 123 572 125
rect 574 123 577 125
rect 569 121 577 123
rect 579 121 584 133
rect 586 131 593 133
rect 618 132 627 137
rect 586 129 589 131
rect 591 129 593 131
rect 586 127 593 129
rect 607 130 614 132
rect 607 128 609 130
rect 611 128 614 130
rect 586 121 592 127
rect 607 126 614 128
rect 524 113 530 119
rect 532 117 539 119
rect 532 115 535 117
rect 537 115 539 117
rect 532 113 539 115
rect 588 119 592 121
rect 609 120 614 126
rect 616 123 627 132
rect 629 123 634 141
rect 636 134 641 141
rect 636 132 643 134
rect 636 130 639 132
rect 641 130 643 132
rect 636 128 643 130
rect 636 123 641 128
rect 616 120 624 123
rect 588 113 594 119
rect 596 117 603 119
rect 596 115 599 117
rect 601 115 603 117
rect 596 113 603 115
rect 650 119 655 125
rect 648 117 655 119
rect 648 115 650 117
rect 652 115 655 117
rect 648 113 655 115
rect 657 123 663 125
rect 657 117 665 123
rect 657 115 660 117
rect 662 115 665 117
rect 657 113 665 115
rect 667 117 675 123
rect 667 115 670 117
rect 672 115 675 117
rect 667 113 675 115
rect 677 121 684 123
rect 677 119 680 121
rect 682 119 684 121
rect 677 113 684 119
rect 4 27 11 33
rect 4 25 6 27
rect 8 25 11 27
rect 4 23 11 25
rect 13 31 21 33
rect 13 29 16 31
rect 18 29 21 31
rect 13 23 21 29
rect 23 31 31 33
rect 23 29 26 31
rect 28 29 31 31
rect 23 23 31 29
rect 25 21 31 23
rect 33 31 40 33
rect 33 29 36 31
rect 38 29 40 31
rect 33 27 40 29
rect 33 21 38 27
rect 85 31 92 33
rect 85 29 87 31
rect 89 29 92 31
rect 85 27 92 29
rect 94 27 100 33
rect 64 23 72 26
rect 47 18 52 23
rect 45 16 52 18
rect 45 14 47 16
rect 49 14 52 16
rect 45 12 52 14
rect 47 5 52 12
rect 54 5 59 23
rect 61 14 72 23
rect 74 20 79 26
rect 96 25 100 27
rect 149 31 156 33
rect 149 29 151 31
rect 153 29 156 31
rect 149 27 156 29
rect 158 27 164 33
rect 74 18 81 20
rect 96 19 102 25
rect 74 16 77 18
rect 79 16 81 18
rect 74 14 81 16
rect 95 17 102 19
rect 95 15 97 17
rect 99 15 102 17
rect 61 9 70 14
rect 95 13 102 15
rect 104 13 109 25
rect 111 23 119 25
rect 111 21 114 23
rect 116 21 119 23
rect 111 13 119 21
rect 121 13 126 25
rect 128 17 136 25
rect 128 15 131 17
rect 133 15 136 17
rect 128 13 136 15
rect 138 23 145 25
rect 138 21 141 23
rect 143 21 145 23
rect 138 19 145 21
rect 160 25 164 27
rect 258 27 264 33
rect 266 31 273 33
rect 266 29 269 31
rect 271 29 273 31
rect 266 27 273 29
rect 258 25 262 27
rect 138 13 143 19
rect 160 19 166 25
rect 159 17 166 19
rect 159 15 161 17
rect 163 15 166 17
rect 159 13 166 15
rect 168 13 173 25
rect 175 23 183 25
rect 175 21 178 23
rect 180 21 183 23
rect 175 13 183 21
rect 185 13 190 25
rect 192 17 200 25
rect 192 15 195 17
rect 197 15 200 17
rect 192 13 200 15
rect 202 23 209 25
rect 202 21 205 23
rect 207 21 209 23
rect 202 19 209 21
rect 213 23 220 25
rect 213 21 215 23
rect 217 21 220 23
rect 213 19 220 21
rect 202 13 207 19
rect 215 13 220 19
rect 222 17 230 25
rect 222 15 225 17
rect 227 15 230 17
rect 222 13 230 15
rect 232 13 237 25
rect 239 23 247 25
rect 239 21 242 23
rect 244 21 247 23
rect 239 13 247 21
rect 249 13 254 25
rect 256 19 262 25
rect 314 32 321 34
rect 314 30 316 32
rect 318 30 321 32
rect 314 28 321 30
rect 323 28 329 34
rect 277 20 285 26
rect 256 17 263 19
rect 256 15 259 17
rect 261 15 263 17
rect 256 13 263 15
rect 276 17 285 20
rect 276 15 278 17
rect 280 15 285 17
rect 61 7 65 9
rect 67 7 70 9
rect 276 10 285 15
rect 276 8 278 10
rect 280 8 285 10
rect 61 5 70 7
rect 276 6 285 8
rect 287 6 292 26
rect 294 18 299 26
rect 325 26 329 28
rect 384 29 389 34
rect 382 27 389 29
rect 325 20 331 26
rect 324 18 331 20
rect 294 16 301 18
rect 294 14 297 16
rect 299 14 301 16
rect 324 16 326 18
rect 328 16 331 18
rect 324 14 331 16
rect 333 14 338 26
rect 340 24 348 26
rect 340 22 343 24
rect 345 22 348 24
rect 340 14 348 22
rect 350 14 355 26
rect 357 18 365 26
rect 357 16 360 18
rect 362 16 365 18
rect 357 14 365 16
rect 367 24 374 26
rect 367 22 370 24
rect 372 22 374 24
rect 367 20 374 22
rect 382 25 384 27
rect 386 25 389 27
rect 382 20 389 25
rect 367 14 372 20
rect 382 18 384 20
rect 386 18 389 20
rect 382 16 389 18
rect 391 27 399 34
rect 423 32 430 34
rect 423 30 425 32
rect 427 30 430 32
rect 391 16 402 27
rect 294 12 301 14
rect 294 6 299 12
rect 393 10 402 16
rect 393 8 395 10
rect 397 8 402 10
rect 393 6 402 8
rect 404 6 409 27
rect 411 19 416 27
rect 423 25 430 30
rect 423 23 425 25
rect 427 23 430 25
rect 423 21 430 23
rect 411 17 418 19
rect 411 15 414 17
rect 416 15 418 17
rect 411 13 418 15
rect 411 6 416 13
rect 425 6 430 21
rect 432 17 440 34
rect 432 15 435 17
rect 437 15 440 17
rect 432 10 440 15
rect 432 8 435 10
rect 437 8 440 10
rect 432 6 440 8
rect 442 25 450 34
rect 442 23 445 25
rect 447 23 450 25
rect 442 18 450 23
rect 442 16 445 18
rect 447 16 450 18
rect 442 6 450 16
rect 452 17 468 34
rect 452 15 457 17
rect 459 15 468 17
rect 452 10 468 15
rect 452 8 457 10
rect 459 9 468 10
rect 470 9 475 34
rect 477 31 482 34
rect 512 32 519 34
rect 477 29 485 31
rect 477 27 480 29
rect 482 27 485 29
rect 477 18 485 27
rect 487 18 498 31
rect 477 9 482 18
rect 489 10 498 18
rect 459 8 466 9
rect 452 6 466 8
rect 489 8 492 10
rect 494 8 498 10
rect 489 6 498 8
rect 500 29 507 31
rect 500 27 503 29
rect 505 27 507 29
rect 500 22 507 27
rect 500 20 503 22
rect 505 20 507 22
rect 512 30 514 32
rect 516 30 519 32
rect 512 25 519 30
rect 512 23 514 25
rect 516 23 519 25
rect 512 21 519 23
rect 500 18 507 20
rect 500 6 505 18
rect 514 6 519 21
rect 521 17 529 34
rect 521 15 524 17
rect 526 15 529 17
rect 521 10 529 15
rect 521 8 524 10
rect 526 8 529 10
rect 521 6 529 8
rect 531 25 539 34
rect 531 23 534 25
rect 536 23 539 25
rect 531 18 539 23
rect 531 16 534 18
rect 536 16 539 18
rect 531 6 539 16
rect 541 17 557 34
rect 541 15 546 17
rect 548 15 557 17
rect 541 10 557 15
rect 541 8 546 10
rect 548 9 557 10
rect 559 9 564 34
rect 566 31 571 34
rect 600 32 607 34
rect 566 29 574 31
rect 566 27 569 29
rect 571 27 574 29
rect 566 18 574 27
rect 576 18 587 31
rect 566 9 571 18
rect 578 10 587 18
rect 548 8 555 9
rect 541 6 555 8
rect 578 8 581 10
rect 583 8 587 10
rect 578 6 587 8
rect 589 29 596 31
rect 589 27 592 29
rect 594 27 596 29
rect 600 30 602 32
rect 604 30 607 32
rect 600 28 607 30
rect 589 22 596 27
rect 602 26 607 28
rect 609 26 615 34
rect 589 20 592 22
rect 594 20 596 22
rect 589 18 596 20
rect 611 22 615 26
rect 664 32 671 34
rect 664 30 666 32
rect 668 30 671 32
rect 664 25 671 30
rect 646 22 651 24
rect 589 6 594 18
rect 611 18 617 22
rect 610 10 617 18
rect 610 8 612 10
rect 614 8 617 10
rect 610 6 617 8
rect 619 6 624 22
rect 626 20 634 22
rect 626 18 629 20
rect 631 18 634 20
rect 626 6 634 18
rect 636 6 641 22
rect 643 10 651 22
rect 643 8 646 10
rect 648 8 651 10
rect 643 6 651 8
rect 653 19 658 24
rect 664 23 666 25
rect 668 23 671 25
rect 664 21 671 23
rect 653 17 660 19
rect 653 15 656 17
rect 658 15 660 17
rect 666 16 671 21
rect 673 17 682 34
rect 673 16 677 17
rect 653 13 660 15
rect 653 6 658 13
rect 675 15 677 16
rect 679 15 682 17
rect 675 13 682 15
<< alu1 >>
rect 0 142 688 146
rect 0 141 418 142
rect 0 139 7 141
rect 9 139 19 141
rect 21 139 301 141
rect 303 139 369 141
rect 371 140 418 141
rect 420 140 534 142
rect 536 140 598 142
rect 600 140 610 142
rect 612 140 651 142
rect 653 140 665 142
rect 667 140 679 142
rect 681 140 688 142
rect 371 139 688 140
rect 0 138 412 139
rect 28 131 41 132
rect 28 129 30 131
rect 32 129 41 131
rect 28 128 41 129
rect 12 123 24 125
rect 12 121 20 123
rect 22 121 24 123
rect 12 119 24 121
rect 20 116 24 119
rect 22 114 24 116
rect 4 107 16 109
rect 4 105 6 107
rect 8 105 13 107
rect 15 105 16 107
rect 4 103 16 105
rect 12 95 16 103
rect 20 102 24 114
rect 20 100 21 102
rect 23 100 24 102
rect 20 98 24 100
rect 22 96 24 98
rect 20 87 24 96
rect 28 107 32 128
rect 83 127 88 133
rect 83 125 84 127
rect 86 125 88 127
rect 28 105 29 107
rect 31 105 32 107
rect 28 95 32 105
rect 83 124 88 125
rect 75 123 88 124
rect 75 121 81 123
rect 83 121 88 123
rect 75 120 88 121
rect 92 128 105 132
rect 181 128 194 132
rect 302 132 306 133
rect 293 128 306 132
rect 92 126 97 128
rect 92 124 94 126
rect 96 124 97 126
rect 181 126 186 128
rect 92 119 97 124
rect 92 117 94 119
rect 96 117 97 119
rect 44 115 56 117
rect 44 113 49 115
rect 51 113 56 115
rect 44 112 56 113
rect 46 111 56 112
rect 46 110 48 111
rect 44 103 48 110
rect 68 107 74 109
rect 68 105 71 107
rect 73 105 74 107
rect 68 100 74 105
rect 68 99 81 100
rect 68 97 69 99
rect 71 97 81 99
rect 68 96 81 97
rect 28 93 33 95
rect 28 91 30 93
rect 32 91 33 93
rect 28 89 33 91
rect 28 87 32 89
rect 92 115 97 117
rect 92 95 96 115
rect 123 115 161 116
rect 123 113 152 115
rect 154 113 161 115
rect 123 112 161 113
rect 123 109 128 112
rect 120 107 128 109
rect 120 105 121 107
rect 123 105 128 107
rect 120 103 128 105
rect 138 107 153 108
rect 138 105 140 107
rect 142 105 147 107
rect 149 105 153 107
rect 138 104 153 105
rect 92 93 93 95
rect 95 93 96 95
rect 92 91 97 93
rect 92 89 94 91
rect 96 89 97 91
rect 92 87 97 89
rect 140 98 144 104
rect 171 123 177 125
rect 171 121 172 123
rect 174 121 177 123
rect 171 116 177 121
rect 171 114 172 116
rect 174 114 177 116
rect 171 112 177 114
rect 140 96 141 98
rect 143 96 144 98
rect 140 87 144 96
rect 173 98 177 112
rect 173 96 174 98
rect 176 96 177 98
rect 173 92 177 96
rect 155 91 177 92
rect 155 89 172 91
rect 174 89 177 91
rect 155 88 177 89
rect 181 124 183 126
rect 185 124 186 126
rect 181 119 186 124
rect 181 117 183 119
rect 185 117 186 119
rect 181 115 186 117
rect 181 113 182 115
rect 184 113 185 115
rect 181 93 185 113
rect 212 112 250 116
rect 212 109 217 112
rect 209 107 217 109
rect 209 105 210 107
rect 212 105 214 107
rect 216 105 217 107
rect 209 103 217 105
rect 227 107 242 108
rect 227 105 229 107
rect 231 105 236 107
rect 238 105 242 107
rect 227 104 242 105
rect 181 91 186 93
rect 229 95 233 104
rect 260 123 266 125
rect 260 121 261 123
rect 263 122 266 123
rect 270 122 274 125
rect 263 121 274 122
rect 260 118 274 121
rect 260 116 266 118
rect 260 114 261 116
rect 263 114 266 116
rect 260 112 266 114
rect 270 116 274 118
rect 270 114 291 116
rect 270 112 275 114
rect 277 112 291 114
rect 262 92 266 112
rect 270 107 291 108
rect 270 105 285 107
rect 287 105 291 107
rect 270 104 291 105
rect 304 126 306 128
rect 369 131 374 133
rect 369 129 370 131
rect 372 129 374 131
rect 302 121 306 126
rect 369 125 374 129
rect 304 119 306 121
rect 270 98 274 104
rect 302 109 306 119
rect 302 107 303 109
rect 305 107 306 109
rect 302 100 306 107
rect 270 96 271 98
rect 273 96 274 98
rect 270 95 274 96
rect 301 98 306 100
rect 301 96 302 98
rect 304 96 306 98
rect 301 94 306 96
rect 314 124 320 125
rect 369 124 370 125
rect 314 122 316 124
rect 318 122 327 124
rect 314 120 327 122
rect 361 123 370 124
rect 372 123 374 125
rect 361 120 374 123
rect 384 132 393 133
rect 384 130 389 132
rect 391 130 393 132
rect 384 129 393 130
rect 181 89 183 91
rect 185 89 186 91
rect 181 87 186 89
rect 244 91 266 92
rect 244 89 261 91
rect 263 89 266 91
rect 244 88 266 89
rect 314 91 318 120
rect 337 110 343 116
rect 328 109 343 110
rect 328 107 330 109
rect 332 107 339 109
rect 341 107 343 109
rect 328 104 343 107
rect 354 107 360 109
rect 354 105 357 107
rect 359 105 360 107
rect 354 101 360 105
rect 354 98 366 101
rect 354 96 360 98
rect 362 96 366 98
rect 354 95 366 96
rect 314 90 320 91
rect 314 88 316 90
rect 318 88 320 90
rect 314 87 320 88
rect 384 112 388 129
rect 415 131 420 133
rect 415 129 416 131
rect 418 129 420 131
rect 415 126 420 129
rect 534 130 539 134
rect 534 128 536 130
rect 538 128 539 130
rect 603 138 607 139
rect 598 131 603 134
rect 598 129 600 131
rect 602 129 603 131
rect 534 126 539 128
rect 598 126 603 129
rect 400 124 404 125
rect 400 122 401 124
rect 403 122 404 124
rect 400 120 404 122
rect 415 124 417 126
rect 419 125 420 126
rect 469 125 475 126
rect 419 124 428 125
rect 415 121 428 124
rect 462 123 471 125
rect 473 123 475 125
rect 462 121 475 123
rect 384 110 385 112
rect 387 110 388 112
rect 392 116 404 120
rect 408 116 412 117
rect 392 115 396 116
rect 392 113 393 115
rect 395 113 396 115
rect 392 111 396 113
rect 408 114 409 116
rect 411 114 412 116
rect 384 107 388 110
rect 408 109 412 114
rect 384 103 396 107
rect 400 106 412 109
rect 400 104 403 106
rect 405 104 412 106
rect 400 103 412 104
rect 392 98 396 103
rect 392 97 401 98
rect 392 95 397 97
rect 399 95 401 97
rect 392 94 401 95
rect 429 108 435 110
rect 429 106 430 108
rect 432 106 435 108
rect 429 102 435 106
rect 423 100 435 102
rect 423 98 429 100
rect 431 98 435 100
rect 423 96 435 98
rect 446 111 452 117
rect 446 110 461 111
rect 446 109 457 110
rect 446 107 452 109
rect 454 108 457 109
rect 459 108 461 110
rect 454 107 461 108
rect 446 105 461 107
rect 471 109 475 121
rect 471 107 472 109
rect 474 107 475 109
rect 471 92 475 107
rect 469 91 475 92
rect 469 89 471 91
rect 473 89 475 91
rect 469 88 475 89
rect 479 125 485 126
rect 534 125 535 126
rect 479 123 481 125
rect 483 123 492 125
rect 479 121 492 123
rect 526 124 535 125
rect 537 124 539 126
rect 526 121 539 124
rect 543 125 549 126
rect 598 125 599 126
rect 543 123 545 125
rect 547 123 556 125
rect 543 121 556 123
rect 590 124 599 125
rect 601 124 603 126
rect 590 121 603 124
rect 607 130 620 133
rect 607 128 609 130
rect 611 129 620 130
rect 479 92 483 121
rect 502 111 508 117
rect 493 110 508 111
rect 493 108 495 110
rect 497 109 508 110
rect 497 108 500 109
rect 493 107 500 108
rect 502 107 508 109
rect 493 105 508 107
rect 519 108 525 110
rect 519 106 522 108
rect 524 106 525 108
rect 519 102 525 106
rect 519 100 531 102
rect 519 98 524 100
rect 526 98 531 100
rect 519 96 531 98
rect 479 91 485 92
rect 479 89 481 91
rect 483 89 485 91
rect 479 88 485 89
rect 543 100 547 121
rect 543 98 544 100
rect 546 98 547 100
rect 543 92 547 98
rect 566 112 572 117
rect 566 111 569 112
rect 557 110 569 111
rect 571 110 572 112
rect 557 108 559 110
rect 561 108 572 110
rect 557 105 572 108
rect 583 108 589 110
rect 583 106 586 108
rect 588 106 589 108
rect 583 102 589 106
rect 583 99 595 102
rect 583 97 592 99
rect 594 97 595 99
rect 583 96 595 97
rect 543 91 549 92
rect 543 89 545 91
rect 547 89 549 91
rect 543 88 549 89
rect 607 112 611 128
rect 607 110 608 112
rect 610 110 611 112
rect 607 96 611 110
rect 631 125 635 126
rect 631 123 632 125
rect 634 123 635 125
rect 631 117 635 123
rect 622 116 635 117
rect 622 114 626 116
rect 628 114 635 116
rect 622 113 635 114
rect 639 109 643 118
rect 630 108 643 109
rect 630 106 636 108
rect 638 106 640 108
rect 642 106 643 108
rect 630 105 643 106
rect 639 104 643 105
rect 648 117 652 126
rect 648 115 650 117
rect 607 94 612 96
rect 607 92 609 94
rect 611 92 612 94
rect 607 88 612 92
rect 648 99 652 115
rect 663 132 676 134
rect 663 130 667 132
rect 669 130 676 132
rect 663 128 676 130
rect 663 125 669 128
rect 663 123 665 125
rect 667 123 669 125
rect 663 121 669 123
rect 680 108 684 110
rect 680 106 681 108
rect 683 106 684 108
rect 648 97 649 99
rect 651 97 652 99
rect 648 94 652 97
rect 648 92 650 94
rect 652 92 660 94
rect 648 88 660 92
rect 680 101 684 106
rect 671 100 684 101
rect 671 98 676 100
rect 678 98 684 100
rect 671 96 684 98
rect 382 82 688 83
rect 0 81 610 82
rect 0 79 7 81
rect 9 79 19 81
rect 21 79 301 81
rect 303 79 387 81
rect 389 79 407 81
rect 409 80 610 81
rect 612 80 638 82
rect 640 80 651 82
rect 653 80 661 82
rect 663 80 688 82
rect 409 79 688 80
rect 0 67 688 79
rect 0 66 279 67
rect 0 64 25 66
rect 27 64 35 66
rect 37 64 48 66
rect 50 64 76 66
rect 78 65 279 66
rect 281 65 299 67
rect 301 65 385 67
rect 387 65 667 67
rect 669 65 679 67
rect 681 65 688 67
rect 78 64 688 65
rect 0 63 305 64
rect 4 48 17 50
rect 4 46 10 48
rect 12 46 17 48
rect 4 45 17 46
rect 4 40 8 45
rect 28 54 40 58
rect 28 52 36 54
rect 38 52 40 54
rect 36 49 40 52
rect 36 47 37 49
rect 39 47 40 49
rect 4 38 5 40
rect 7 38 8 40
rect 4 36 8 38
rect 19 23 25 25
rect 19 21 21 23
rect 23 21 25 23
rect 19 18 25 21
rect 12 16 25 18
rect 12 14 19 16
rect 21 14 25 16
rect 12 12 25 14
rect 36 31 40 47
rect 76 54 81 58
rect 76 52 77 54
rect 79 52 81 54
rect 76 50 81 52
rect 38 29 40 31
rect 36 20 40 29
rect 45 41 49 42
rect 45 40 58 41
rect 45 38 46 40
rect 48 38 50 40
rect 52 38 58 40
rect 45 37 58 38
rect 45 28 49 37
rect 53 32 66 33
rect 53 30 60 32
rect 62 30 66 32
rect 53 29 66 30
rect 53 23 57 29
rect 53 21 54 23
rect 56 21 57 23
rect 53 20 57 21
rect 77 36 81 50
rect 77 34 78 36
rect 80 34 81 36
rect 77 18 81 34
rect 139 57 145 58
rect 139 55 141 57
rect 143 55 145 57
rect 139 54 145 55
rect 93 49 105 50
rect 93 47 94 49
rect 96 47 105 49
rect 93 44 105 47
rect 99 40 105 44
rect 99 38 100 40
rect 102 38 105 40
rect 99 36 105 38
rect 116 38 131 41
rect 116 36 127 38
rect 129 36 131 38
rect 116 34 117 36
rect 119 35 131 36
rect 119 34 122 35
rect 116 29 122 34
rect 141 48 145 54
rect 141 46 142 48
rect 144 46 145 48
rect 141 25 145 46
rect 203 57 209 58
rect 203 55 205 57
rect 207 55 209 57
rect 203 54 209 55
rect 157 48 169 50
rect 157 46 162 48
rect 164 46 169 48
rect 157 44 169 46
rect 163 40 169 44
rect 163 38 164 40
rect 166 38 169 40
rect 163 36 169 38
rect 180 39 195 41
rect 180 37 186 39
rect 188 38 195 39
rect 188 37 191 38
rect 180 36 191 37
rect 193 36 195 38
rect 180 35 195 36
rect 180 29 186 35
rect 205 25 209 54
rect 68 16 77 17
rect 79 16 81 18
rect 68 13 81 16
rect 85 22 98 25
rect 85 20 87 22
rect 89 21 98 22
rect 132 23 145 25
rect 132 21 141 23
rect 143 21 145 23
rect 89 20 90 21
rect 139 20 145 21
rect 149 22 162 25
rect 149 20 151 22
rect 153 21 162 22
rect 196 23 209 25
rect 196 21 205 23
rect 207 21 209 23
rect 153 20 154 21
rect 203 20 209 21
rect 213 57 219 58
rect 213 55 215 57
rect 217 55 219 57
rect 213 54 219 55
rect 213 39 217 54
rect 213 37 214 39
rect 216 37 217 39
rect 213 25 217 37
rect 227 39 242 41
rect 227 38 234 39
rect 227 36 229 38
rect 231 37 234 38
rect 236 37 242 39
rect 231 36 242 37
rect 227 35 242 36
rect 236 29 242 35
rect 253 48 265 50
rect 253 46 257 48
rect 259 46 265 48
rect 253 44 265 46
rect 253 40 259 44
rect 253 38 256 40
rect 258 38 259 40
rect 253 36 259 38
rect 287 51 296 52
rect 287 49 289 51
rect 291 49 296 51
rect 287 48 296 49
rect 292 43 296 48
rect 276 42 288 43
rect 276 40 283 42
rect 285 40 288 42
rect 276 37 288 40
rect 292 39 304 43
rect 276 32 280 37
rect 300 36 304 39
rect 276 30 277 32
rect 279 30 280 32
rect 292 33 296 35
rect 292 31 293 33
rect 295 31 296 33
rect 292 30 296 31
rect 276 29 280 30
rect 284 26 296 30
rect 300 34 301 36
rect 303 34 304 36
rect 213 23 226 25
rect 213 21 215 23
rect 217 21 226 23
rect 260 22 273 25
rect 260 21 269 22
rect 213 20 219 21
rect 268 20 269 21
rect 271 20 273 22
rect 284 24 288 26
rect 284 22 285 24
rect 287 22 288 24
rect 284 21 288 22
rect 85 17 90 20
rect 149 18 154 20
rect 85 15 86 17
rect 88 15 90 17
rect 85 12 90 15
rect 81 7 85 8
rect 149 16 150 18
rect 152 16 154 18
rect 149 12 154 16
rect 268 17 273 20
rect 268 15 270 17
rect 272 15 273 17
rect 268 13 273 15
rect 300 17 304 34
rect 368 58 378 59
rect 368 56 370 58
rect 372 56 375 58
rect 377 56 378 58
rect 368 55 378 56
rect 370 53 378 55
rect 422 57 444 58
rect 422 55 425 57
rect 427 55 444 57
rect 422 54 444 55
rect 502 57 507 59
rect 502 55 503 57
rect 505 55 507 57
rect 322 50 334 51
rect 322 48 326 50
rect 328 48 334 50
rect 322 45 334 48
rect 328 41 334 45
rect 328 39 329 41
rect 331 39 334 41
rect 328 37 334 39
rect 345 39 360 42
rect 345 37 347 39
rect 349 37 356 39
rect 358 37 360 39
rect 345 36 360 37
rect 345 30 351 36
rect 370 26 374 53
rect 295 16 304 17
rect 295 14 297 16
rect 299 14 304 16
rect 295 13 304 14
rect 314 23 327 26
rect 314 21 316 23
rect 318 22 327 23
rect 361 24 374 26
rect 361 22 370 24
rect 372 22 374 24
rect 318 21 319 22
rect 368 21 374 22
rect 382 50 387 52
rect 382 48 384 50
rect 386 48 387 50
rect 382 46 387 48
rect 414 50 418 51
rect 414 48 415 50
rect 417 48 418 50
rect 382 39 386 46
rect 382 37 383 39
rect 385 37 386 39
rect 382 27 386 37
rect 414 42 418 48
rect 382 25 384 27
rect 314 17 319 21
rect 382 20 386 25
rect 314 15 316 17
rect 318 15 319 17
rect 314 13 319 15
rect 382 18 384 20
rect 397 41 418 42
rect 397 39 401 41
rect 403 39 418 41
rect 397 38 418 39
rect 422 34 426 54
rect 397 32 411 34
rect 413 32 418 34
rect 397 30 418 32
rect 414 28 418 30
rect 422 32 428 34
rect 422 30 425 32
rect 427 30 428 32
rect 422 28 428 30
rect 414 25 428 28
rect 414 24 425 25
rect 414 21 418 24
rect 422 23 425 24
rect 427 23 428 25
rect 422 21 428 23
rect 455 42 459 51
rect 502 53 507 55
rect 446 41 461 42
rect 446 39 450 41
rect 452 39 457 41
rect 459 39 461 41
rect 446 38 461 39
rect 471 41 479 43
rect 471 39 472 41
rect 474 39 476 41
rect 478 39 479 41
rect 471 37 479 39
rect 471 34 476 37
rect 438 30 476 34
rect 503 33 507 53
rect 503 31 504 33
rect 506 31 507 33
rect 502 29 507 31
rect 502 27 503 29
rect 505 27 507 29
rect 502 22 507 27
rect 502 20 503 22
rect 505 20 507 22
rect 511 57 533 58
rect 511 55 514 57
rect 516 55 533 57
rect 511 54 533 55
rect 511 50 515 54
rect 511 48 512 50
rect 514 48 515 50
rect 511 34 515 48
rect 544 50 548 59
rect 544 48 545 50
rect 547 48 548 50
rect 511 32 517 34
rect 511 30 514 32
rect 516 30 517 32
rect 511 25 517 30
rect 511 23 514 25
rect 516 23 517 25
rect 511 21 517 23
rect 544 42 548 48
rect 591 57 596 59
rect 591 55 592 57
rect 594 55 596 57
rect 591 53 596 55
rect 592 51 593 53
rect 595 51 596 53
rect 535 41 550 42
rect 535 39 539 41
rect 541 39 546 41
rect 548 39 550 41
rect 535 38 550 39
rect 560 41 568 43
rect 560 39 565 41
rect 567 39 568 41
rect 560 37 568 39
rect 560 34 565 37
rect 527 33 565 34
rect 527 31 534 33
rect 536 31 565 33
rect 527 30 565 31
rect 592 31 596 51
rect 591 29 596 31
rect 656 57 660 59
rect 655 55 660 57
rect 655 53 656 55
rect 658 53 660 55
rect 655 51 660 53
rect 607 49 620 50
rect 607 47 617 49
rect 619 47 620 49
rect 607 46 620 47
rect 614 41 620 46
rect 614 39 615 41
rect 617 39 620 41
rect 614 37 620 39
rect 640 36 644 43
rect 640 35 642 36
rect 632 34 642 35
rect 632 33 644 34
rect 632 31 637 33
rect 639 31 644 33
rect 632 29 644 31
rect 591 27 592 29
rect 594 27 596 29
rect 591 22 596 27
rect 502 18 507 20
rect 591 20 592 22
rect 594 20 596 22
rect 591 18 596 20
rect 382 14 395 18
rect 382 13 386 14
rect 494 14 507 18
rect 583 14 596 18
rect 600 25 613 26
rect 600 23 602 25
rect 604 23 613 25
rect 600 22 613 23
rect 600 21 605 22
rect 656 41 660 51
rect 656 39 657 41
rect 659 39 660 41
rect 600 19 602 21
rect 604 19 605 21
rect 600 13 605 19
rect 656 18 660 39
rect 664 50 668 59
rect 664 48 666 50
rect 664 46 668 48
rect 664 44 665 46
rect 667 44 668 46
rect 664 32 668 44
rect 672 43 676 51
rect 672 41 684 43
rect 672 39 673 41
rect 675 39 680 41
rect 682 39 684 41
rect 672 37 684 39
rect 664 30 666 32
rect 664 27 668 30
rect 664 25 676 27
rect 664 23 666 25
rect 668 23 676 25
rect 664 21 676 23
rect 647 17 660 18
rect 647 15 656 17
rect 658 15 660 17
rect 647 14 660 15
rect 276 7 688 8
rect 0 6 317 7
rect 0 4 7 6
rect 9 4 21 6
rect 23 4 35 6
rect 37 4 76 6
rect 78 4 88 6
rect 90 4 152 6
rect 154 4 268 6
rect 270 5 317 6
rect 319 5 385 7
rect 387 5 667 7
rect 669 5 679 7
rect 681 5 688 7
rect 270 4 688 5
rect 0 0 688 4
<< alu2 >>
rect 524 135 547 139
rect 369 131 374 133
rect 524 132 528 135
rect 369 129 370 131
rect 372 129 374 131
rect 83 124 88 125
rect 77 123 84 124
rect 77 121 81 123
rect 83 122 84 123
rect 86 122 88 124
rect 83 121 88 122
rect 77 120 88 121
rect 4 115 52 116
rect 4 113 49 115
rect 51 113 52 115
rect 4 112 52 113
rect 151 115 185 116
rect 151 113 152 115
rect 154 113 182 115
rect 184 113 185 115
rect 151 112 185 113
rect 4 107 9 112
rect 302 109 343 110
rect 4 105 6 107
rect 8 105 9 107
rect 4 42 9 105
rect 28 107 217 108
rect 28 105 29 107
rect 31 105 214 107
rect 216 105 217 107
rect 302 107 303 109
rect 305 107 339 109
rect 341 107 343 109
rect 302 106 343 107
rect 28 104 217 105
rect 20 102 24 103
rect 20 100 21 102
rect 23 100 24 102
rect 20 99 72 100
rect 20 97 69 99
rect 71 97 72 99
rect 20 96 72 97
rect 140 98 144 100
rect 140 96 141 98
rect 143 96 144 98
rect 92 95 96 96
rect 92 93 93 95
rect 95 93 96 95
rect 92 82 96 93
rect 140 91 144 96
rect 173 98 364 99
rect 173 96 174 98
rect 176 96 178 98
rect 180 96 271 98
rect 273 96 360 98
rect 362 96 364 98
rect 173 95 364 96
rect 140 89 141 91
rect 143 89 265 91
rect 140 87 265 89
rect 92 78 232 82
rect 36 49 97 50
rect 36 47 37 49
rect 39 47 94 49
rect 96 47 97 49
rect 36 46 97 47
rect 141 48 169 50
rect 141 46 142 48
rect 144 46 162 48
rect 164 46 169 48
rect 141 44 169 46
rect 4 40 49 42
rect 227 41 232 78
rect 259 50 265 87
rect 369 80 374 129
rect 400 131 528 132
rect 543 132 547 135
rect 543 131 603 132
rect 400 129 416 131
rect 418 129 528 131
rect 400 128 528 129
rect 533 130 539 131
rect 533 128 536 130
rect 538 128 539 130
rect 543 129 600 131
rect 602 129 603 131
rect 543 128 603 129
rect 400 124 404 128
rect 533 124 539 128
rect 400 122 401 124
rect 403 122 404 124
rect 400 121 404 122
rect 408 120 539 124
rect 630 125 669 126
rect 630 123 632 125
rect 634 123 665 125
rect 667 123 669 125
rect 630 122 669 123
rect 408 116 412 120
rect 630 117 635 122
rect 300 75 374 80
rect 384 112 388 115
rect 408 114 409 116
rect 411 114 412 116
rect 408 112 412 114
rect 622 116 635 117
rect 622 114 623 116
rect 625 114 635 116
rect 622 113 635 114
rect 567 112 611 113
rect 384 110 385 112
rect 387 110 388 112
rect 253 48 271 50
rect 253 46 257 48
rect 259 46 271 48
rect 253 44 271 46
rect 4 38 5 40
rect 7 38 46 40
rect 48 38 49 40
rect 4 36 49 38
rect 180 39 217 41
rect 180 37 186 39
rect 188 37 214 39
rect 216 37 217 39
rect 77 36 121 37
rect 77 34 78 36
rect 80 34 117 36
rect 119 34 121 36
rect 180 35 217 37
rect 227 39 239 41
rect 227 37 234 39
rect 236 37 239 39
rect 227 35 239 37
rect 300 36 304 75
rect 384 70 388 110
rect 449 109 461 111
rect 449 107 452 109
rect 454 107 461 109
rect 449 105 461 107
rect 471 109 508 111
rect 567 110 569 112
rect 571 110 608 112
rect 610 110 611 112
rect 567 109 611 110
rect 471 107 472 109
rect 474 107 500 109
rect 502 107 508 109
rect 471 105 508 107
rect 639 108 684 110
rect 639 106 640 108
rect 642 106 681 108
rect 683 106 684 108
rect 417 100 435 102
rect 417 98 429 100
rect 431 98 435 100
rect 417 96 435 98
rect 300 34 301 36
rect 303 34 304 36
rect 77 33 121 34
rect 53 32 66 33
rect 53 30 63 32
rect 65 30 66 32
rect 53 29 66 30
rect 276 32 280 34
rect 276 30 277 32
rect 279 30 280 32
rect 300 31 304 34
rect 314 65 388 70
rect 53 24 58 29
rect 276 26 280 30
rect 19 23 58 24
rect 19 21 21 23
rect 23 21 54 23
rect 56 21 58 23
rect 19 20 58 21
rect 149 22 280 26
rect 284 24 288 25
rect 284 22 285 24
rect 287 22 288 24
rect 149 18 155 22
rect 284 18 288 22
rect 85 17 145 18
rect 85 15 86 17
rect 88 15 145 17
rect 149 16 150 18
rect 152 16 155 18
rect 149 15 155 16
rect 160 17 288 18
rect 160 15 270 17
rect 272 15 288 17
rect 85 14 145 15
rect 141 11 145 14
rect 160 14 288 15
rect 314 17 319 65
rect 370 60 379 61
rect 370 58 371 60
rect 373 58 379 60
rect 370 56 375 58
rect 377 56 379 58
rect 370 55 379 56
rect 423 59 429 96
rect 456 68 461 105
rect 639 104 684 106
rect 519 100 547 102
rect 519 98 524 100
rect 526 98 544 100
rect 546 98 547 100
rect 519 96 547 98
rect 591 99 652 100
rect 591 97 592 99
rect 594 97 649 99
rect 651 97 652 99
rect 591 96 652 97
rect 456 64 596 68
rect 423 55 548 59
rect 544 53 548 55
rect 544 51 545 53
rect 547 51 548 53
rect 324 50 515 51
rect 324 48 326 50
rect 328 48 415 50
rect 417 48 508 50
rect 510 48 512 50
rect 514 48 515 50
rect 324 47 515 48
rect 544 50 548 51
rect 592 53 596 64
rect 592 51 593 53
rect 595 51 596 53
rect 592 50 596 51
rect 544 48 545 50
rect 547 48 548 50
rect 544 46 548 48
rect 616 49 668 50
rect 616 47 617 49
rect 619 47 668 49
rect 616 46 668 47
rect 664 44 665 46
rect 667 44 668 46
rect 664 43 668 44
rect 471 41 660 42
rect 345 39 386 40
rect 345 37 347 39
rect 349 37 383 39
rect 385 37 386 39
rect 471 39 472 41
rect 474 39 657 41
rect 659 39 660 41
rect 471 38 660 39
rect 679 41 684 104
rect 679 39 680 41
rect 682 39 684 41
rect 345 36 386 37
rect 679 34 684 39
rect 503 33 537 34
rect 503 31 504 33
rect 506 31 534 33
rect 536 31 537 33
rect 503 30 537 31
rect 636 33 684 34
rect 636 31 637 33
rect 639 31 684 33
rect 636 30 684 31
rect 314 15 316 17
rect 318 15 319 17
rect 160 11 164 14
rect 314 13 319 15
rect 600 25 605 26
rect 600 23 602 25
rect 604 23 605 25
rect 600 16 605 23
rect 600 14 601 16
rect 603 14 605 16
rect 600 13 605 14
rect 141 7 164 11
<< alu3 >>
rect 83 131 88 133
rect 83 129 84 131
rect 86 129 88 131
rect 83 124 88 129
rect 79 122 84 124
rect 86 122 88 124
rect 79 120 88 122
rect 622 116 626 117
rect 622 114 623 116
rect 625 114 626 116
rect 140 94 144 102
rect 140 92 141 94
rect 143 92 144 94
rect 140 91 144 92
rect 140 89 141 91
rect 143 89 144 91
rect 140 87 144 89
rect 177 98 181 99
rect 177 96 178 98
rect 180 96 181 98
rect 177 75 181 96
rect 622 75 626 114
rect 62 71 181 75
rect 507 71 626 75
rect 62 32 66 71
rect 370 60 376 61
rect 370 58 371 60
rect 373 58 376 60
rect 370 57 376 58
rect 370 55 371 57
rect 373 55 376 57
rect 370 53 376 55
rect 507 50 511 71
rect 507 48 508 50
rect 510 48 511 50
rect 507 47 511 48
rect 544 53 548 59
rect 544 51 545 53
rect 547 51 548 53
rect 62 30 63 32
rect 65 30 66 32
rect 62 29 66 30
rect 544 17 548 51
rect 544 16 605 17
rect 544 14 601 16
rect 603 14 605 16
rect 544 12 545 14
rect 547 13 605 14
rect 547 12 550 13
rect 544 10 550 12
<< alu4 >>
rect 83 131 88 133
rect 83 129 84 131
rect 86 129 88 131
rect 36 45 40 49
rect 83 17 88 129
rect 648 97 652 101
rect 140 94 144 97
rect 140 92 141 94
rect 143 92 144 94
rect 140 73 144 92
rect 140 68 374 73
rect 370 57 374 68
rect 370 55 371 57
rect 373 55 374 57
rect 370 51 374 55
rect 83 14 550 17
rect 83 12 545 14
rect 547 12 550 14
rect 83 10 550 12
<< ptie >>
rect 5 81 23 83
rect 5 79 7 81
rect 9 79 19 81
rect 21 79 23 81
rect 5 77 23 79
rect 299 81 305 83
rect 299 79 301 81
rect 303 79 305 81
rect 299 77 305 79
rect 385 81 411 83
rect 385 79 387 81
rect 389 79 407 81
rect 409 79 411 81
rect 385 77 411 79
rect 608 82 642 84
rect 608 80 610 82
rect 612 80 638 82
rect 640 80 642 82
rect 608 78 642 80
rect 649 82 655 84
rect 649 80 651 82
rect 653 80 655 82
rect 649 78 655 80
rect 33 66 39 68
rect 33 64 35 66
rect 37 64 39 66
rect 33 62 39 64
rect 46 66 80 68
rect 46 64 48 66
rect 50 64 76 66
rect 78 64 80 66
rect 46 62 80 64
rect 277 67 303 69
rect 277 65 279 67
rect 281 65 299 67
rect 301 65 303 67
rect 277 63 303 65
rect 383 67 389 69
rect 383 65 385 67
rect 387 65 389 67
rect 383 63 389 65
rect 665 67 683 69
rect 665 65 667 67
rect 669 65 679 67
rect 681 65 683 67
rect 665 63 683 65
<< ntie >>
rect 5 141 23 143
rect 5 139 7 141
rect 9 139 19 141
rect 21 139 23 141
rect 5 137 23 139
rect 299 141 305 143
rect 299 139 301 141
rect 303 139 305 141
rect 299 137 305 139
rect 367 141 373 143
rect 367 139 369 141
rect 371 139 373 141
rect 416 142 422 144
rect 416 140 418 142
rect 420 140 422 142
rect 367 137 373 139
rect 416 138 422 140
rect 532 142 538 144
rect 532 140 534 142
rect 536 140 538 142
rect 532 138 538 140
rect 596 142 602 144
rect 596 140 598 142
rect 600 140 602 142
rect 596 138 602 140
rect 608 142 614 144
rect 608 140 610 142
rect 612 140 614 142
rect 649 142 683 144
rect 608 138 614 140
rect 649 140 651 142
rect 653 140 665 142
rect 667 140 679 142
rect 681 140 683 142
rect 649 138 683 140
rect 5 6 39 8
rect 5 4 7 6
rect 9 4 21 6
rect 23 4 35 6
rect 37 4 39 6
rect 74 6 80 8
rect 5 2 39 4
rect 74 4 76 6
rect 78 4 80 6
rect 74 2 80 4
rect 86 6 92 8
rect 86 4 88 6
rect 90 4 92 6
rect 86 2 92 4
rect 150 6 156 8
rect 150 4 152 6
rect 154 4 156 6
rect 150 2 156 4
rect 266 6 272 8
rect 315 7 321 9
rect 266 4 268 6
rect 270 4 272 6
rect 266 2 272 4
rect 315 5 317 7
rect 319 5 321 7
rect 315 3 321 5
rect 383 7 389 9
rect 383 5 385 7
rect 387 5 389 7
rect 383 3 389 5
rect 665 7 683 9
rect 665 5 667 7
rect 669 5 679 7
rect 681 5 683 7
rect 665 3 683 5
<< nmos >>
rect 15 91 17 100
rect 35 86 37 95
rect 45 86 47 94
rect 52 86 54 94
rect 62 86 64 94
rect 69 86 71 94
rect 79 88 81 94
rect 99 80 101 93
rect 109 83 111 93
rect 119 86 121 100
rect 129 86 131 100
rect 149 80 151 100
rect 156 80 158 100
rect 167 80 169 94
rect 188 80 190 93
rect 198 83 200 93
rect 208 86 210 100
rect 218 86 220 100
rect 238 80 240 100
rect 245 80 247 100
rect 277 94 279 100
rect 287 94 289 100
rect 256 80 258 94
rect 297 91 299 100
rect 392 93 394 99
rect 402 93 404 99
rect 321 86 323 92
rect 331 86 333 92
rect 338 86 340 92
rect 348 86 350 92
rect 355 86 357 92
rect 365 86 367 92
rect 422 87 424 93
rect 432 87 434 93
rect 439 87 441 93
rect 449 87 451 93
rect 456 87 458 93
rect 466 87 468 93
rect 486 87 488 93
rect 496 87 498 93
rect 503 87 505 93
rect 513 87 515 93
rect 520 87 522 93
rect 530 87 532 93
rect 550 87 552 93
rect 560 87 562 93
rect 567 87 569 93
rect 577 87 579 93
rect 584 87 586 93
rect 594 87 596 93
rect 614 90 616 96
rect 624 90 626 96
rect 634 90 636 96
rect 655 90 657 96
rect 667 84 669 93
rect 674 84 676 93
rect 12 53 14 62
rect 19 53 21 62
rect 31 50 33 56
rect 52 50 54 56
rect 62 50 64 56
rect 72 50 74 56
rect 92 53 94 59
rect 102 53 104 59
rect 109 53 111 59
rect 119 53 121 59
rect 126 53 128 59
rect 136 53 138 59
rect 156 53 158 59
rect 166 53 168 59
rect 173 53 175 59
rect 183 53 185 59
rect 190 53 192 59
rect 200 53 202 59
rect 220 53 222 59
rect 230 53 232 59
rect 237 53 239 59
rect 247 53 249 59
rect 254 53 256 59
rect 264 53 266 59
rect 321 54 323 60
rect 331 54 333 60
rect 338 54 340 60
rect 348 54 350 60
rect 355 54 357 60
rect 365 54 367 60
rect 284 47 286 53
rect 294 47 296 53
rect 389 46 391 55
rect 430 52 432 66
rect 399 46 401 52
rect 409 46 411 52
rect 441 46 443 66
rect 448 46 450 66
rect 468 46 470 60
rect 478 46 480 60
rect 488 53 490 63
rect 498 53 500 66
rect 519 52 521 66
rect 530 46 532 66
rect 537 46 539 66
rect 557 46 559 60
rect 567 46 569 60
rect 577 53 579 63
rect 587 53 589 66
rect 607 52 609 58
rect 617 52 619 60
rect 624 52 626 60
rect 634 52 636 60
rect 641 52 643 60
rect 651 51 653 60
rect 671 46 673 55
<< pmos >>
rect 15 112 17 130
rect 35 122 37 140
rect 45 124 47 140
rect 52 124 54 140
rect 62 124 64 140
rect 69 124 71 140
rect 79 112 81 120
rect 99 115 101 140
rect 112 115 114 128
rect 122 112 124 137
rect 129 112 131 137
rect 147 112 149 140
rect 157 112 159 140
rect 167 112 169 140
rect 188 115 190 140
rect 201 115 203 128
rect 211 112 213 137
rect 218 112 220 137
rect 236 112 238 140
rect 246 112 248 140
rect 256 112 258 140
rect 277 119 279 140
rect 284 119 286 140
rect 297 112 299 130
rect 321 120 323 132
rect 331 120 333 132
rect 338 120 340 132
rect 348 120 350 132
rect 355 120 357 132
rect 394 120 396 140
rect 401 120 403 140
rect 365 112 367 118
rect 432 121 434 133
rect 439 121 441 133
rect 449 121 451 133
rect 456 121 458 133
rect 466 121 468 133
rect 486 121 488 133
rect 496 121 498 133
rect 503 121 505 133
rect 513 121 515 133
rect 520 121 522 133
rect 422 113 424 119
rect 550 121 552 133
rect 560 121 562 133
rect 567 121 569 133
rect 577 121 579 133
rect 584 121 586 133
rect 530 113 532 119
rect 614 120 616 132
rect 627 123 629 141
rect 634 123 636 141
rect 594 113 596 119
rect 655 113 657 125
rect 665 113 667 123
rect 675 113 677 123
rect 11 23 13 33
rect 21 23 23 33
rect 31 21 33 33
rect 92 27 94 33
rect 52 5 54 23
rect 59 5 61 23
rect 72 14 74 26
rect 156 27 158 33
rect 102 13 104 25
rect 109 13 111 25
rect 119 13 121 25
rect 126 13 128 25
rect 136 13 138 25
rect 264 27 266 33
rect 166 13 168 25
rect 173 13 175 25
rect 183 13 185 25
rect 190 13 192 25
rect 200 13 202 25
rect 220 13 222 25
rect 230 13 232 25
rect 237 13 239 25
rect 247 13 249 25
rect 254 13 256 25
rect 321 28 323 34
rect 285 6 287 26
rect 292 6 294 26
rect 331 14 333 26
rect 338 14 340 26
rect 348 14 350 26
rect 355 14 357 26
rect 365 14 367 26
rect 389 16 391 34
rect 402 6 404 27
rect 409 6 411 27
rect 430 6 432 34
rect 440 6 442 34
rect 450 6 452 34
rect 468 9 470 34
rect 475 9 477 34
rect 485 18 487 31
rect 498 6 500 31
rect 519 6 521 34
rect 529 6 531 34
rect 539 6 541 34
rect 557 9 559 34
rect 564 9 566 34
rect 574 18 576 31
rect 587 6 589 31
rect 607 26 609 34
rect 617 6 619 22
rect 624 6 626 22
rect 634 6 636 22
rect 641 6 643 22
rect 651 6 653 24
rect 671 16 673 34
<< polyct0 >>
rect 61 115 63 117
rect 36 100 38 102
rect 54 99 56 101
rect 107 108 109 110
rect 101 98 103 100
rect 157 105 159 107
rect 167 105 169 107
rect 196 108 198 110
rect 190 98 192 100
rect 246 105 248 107
rect 256 105 258 107
rect 295 105 297 107
rect 347 113 349 115
rect 322 97 324 99
rect 340 97 342 99
rect 440 114 442 116
rect 447 98 449 100
rect 512 114 514 116
rect 465 98 467 100
rect 487 98 489 100
rect 505 98 507 100
rect 576 114 578 116
rect 551 98 553 100
rect 569 98 571 100
rect 616 107 618 109
rect 657 106 659 108
rect 29 38 31 40
rect 70 37 72 39
rect 117 46 119 48
rect 135 46 137 48
rect 110 30 112 32
rect 181 46 183 48
rect 199 46 201 48
rect 221 46 223 48
rect 174 30 176 32
rect 239 46 241 48
rect 246 30 248 32
rect 346 47 348 49
rect 364 47 366 49
rect 339 31 341 33
rect 391 39 393 41
rect 430 39 432 41
rect 440 39 442 41
rect 496 46 498 48
rect 490 36 492 38
rect 519 39 521 41
rect 529 39 531 41
rect 585 46 587 48
rect 579 36 581 38
rect 632 45 634 47
rect 650 44 652 46
rect 625 29 627 31
<< polyct1 >>
rect 84 125 86 127
rect 13 105 15 107
rect 44 110 46 112
rect 71 105 73 107
rect 121 105 123 107
rect 140 105 142 107
rect 147 105 149 107
rect 275 112 277 114
rect 210 105 212 107
rect 229 105 231 107
rect 236 105 238 107
rect 370 123 372 125
rect 285 105 287 107
rect 330 107 332 109
rect 417 124 419 126
rect 393 113 395 115
rect 357 105 359 107
rect 535 124 537 126
rect 403 104 405 106
rect 430 106 432 108
rect 457 108 459 110
rect 495 108 497 110
rect 599 124 601 126
rect 522 106 524 108
rect 559 108 561 110
rect 667 130 669 132
rect 586 106 588 108
rect 626 114 628 116
rect 636 106 638 108
rect 676 98 678 100
rect 10 46 12 48
rect 50 38 52 40
rect 60 30 62 32
rect 100 38 102 40
rect 19 14 21 16
rect 127 36 129 38
rect 164 38 166 40
rect 87 20 89 22
rect 191 36 193 38
rect 229 36 231 38
rect 256 38 258 40
rect 283 40 285 42
rect 151 20 153 22
rect 329 39 331 41
rect 293 31 295 33
rect 269 20 271 22
rect 356 37 358 39
rect 401 39 403 41
rect 316 21 318 23
rect 450 39 452 41
rect 457 39 459 41
rect 476 39 478 41
rect 411 32 413 34
rect 539 39 541 41
rect 546 39 548 41
rect 565 39 567 41
rect 615 39 617 41
rect 642 34 644 36
rect 673 39 675 41
rect 602 19 604 21
<< ndifct0 >>
rect 6 93 8 95
rect 40 88 42 90
rect 57 88 59 90
rect 74 90 76 92
rect 84 90 86 92
rect 104 85 106 87
rect 114 88 116 90
rect 124 96 126 98
rect 134 96 136 98
rect 134 89 136 91
rect 144 89 146 91
rect 161 82 163 84
rect 193 85 195 87
rect 203 88 205 90
rect 213 96 215 98
rect 223 96 225 98
rect 223 89 225 91
rect 233 89 235 91
rect 282 96 284 98
rect 250 82 252 84
rect 386 95 388 97
rect 407 95 409 97
rect 272 83 274 85
rect 326 88 328 90
rect 343 88 345 90
rect 360 88 362 90
rect 370 88 372 90
rect 417 89 419 91
rect 427 89 429 91
rect 444 89 446 91
rect 461 89 463 91
rect 491 89 493 91
rect 508 89 510 91
rect 525 89 527 91
rect 535 89 537 91
rect 555 89 557 91
rect 572 89 574 91
rect 589 89 591 91
rect 599 89 601 91
rect 619 92 621 94
rect 629 92 631 94
rect 639 92 641 94
rect 291 83 293 85
rect 679 89 681 91
rect 7 55 9 57
rect 395 61 397 63
rect 47 52 49 54
rect 57 52 59 54
rect 67 52 69 54
rect 87 55 89 57
rect 97 55 99 57
rect 114 55 116 57
rect 131 55 133 57
rect 151 55 153 57
rect 161 55 163 57
rect 178 55 180 57
rect 195 55 197 57
rect 225 55 227 57
rect 242 55 244 57
rect 259 55 261 57
rect 269 55 271 57
rect 316 56 318 58
rect 326 56 328 58
rect 343 56 345 58
rect 360 56 362 58
rect 414 61 416 63
rect 279 49 281 51
rect 300 49 302 51
rect 436 62 438 64
rect 404 48 406 50
rect 453 55 455 57
rect 463 55 465 57
rect 463 48 465 50
rect 473 48 475 50
rect 483 56 485 58
rect 493 59 495 61
rect 525 62 527 64
rect 542 55 544 57
rect 552 55 554 57
rect 552 48 554 50
rect 562 48 564 50
rect 572 56 574 58
rect 582 59 584 61
rect 602 54 604 56
rect 612 54 614 56
rect 629 56 631 58
rect 646 56 648 58
rect 680 51 682 53
<< ndifct1 >>
rect 20 96 22 98
rect 30 91 32 93
rect 94 89 96 91
rect 172 89 174 91
rect 183 89 185 91
rect 261 89 263 91
rect 302 96 304 98
rect 397 95 399 97
rect 316 88 318 90
rect 471 89 473 91
rect 481 89 483 91
rect 545 89 547 91
rect 609 92 611 94
rect 650 92 652 94
rect 661 80 663 82
rect 25 64 27 66
rect 36 52 38 54
rect 77 52 79 54
rect 141 55 143 57
rect 205 55 207 57
rect 215 55 217 57
rect 370 56 372 58
rect 289 49 291 51
rect 384 48 386 50
rect 425 55 427 57
rect 503 55 505 57
rect 514 55 516 57
rect 592 55 594 57
rect 656 53 658 55
rect 666 48 668 50
<< ntiect1 >>
rect 7 139 9 141
rect 19 139 21 141
rect 301 139 303 141
rect 369 139 371 141
rect 418 140 420 142
rect 534 140 536 142
rect 598 140 600 142
rect 610 140 612 142
rect 651 140 653 142
rect 665 140 667 142
rect 679 140 681 142
rect 7 4 9 6
rect 21 4 23 6
rect 35 4 37 6
rect 76 4 78 6
rect 88 4 90 6
rect 152 4 154 6
rect 268 4 270 6
rect 317 5 319 7
rect 385 5 387 7
rect 667 5 669 7
rect 679 5 681 7
<< ptiect1 >>
rect 7 79 9 81
rect 19 79 21 81
rect 301 79 303 81
rect 387 79 389 81
rect 407 79 409 81
rect 610 80 612 82
rect 638 80 640 82
rect 651 80 653 82
rect 35 64 37 66
rect 48 64 50 66
rect 76 64 78 66
rect 279 65 281 67
rect 299 65 301 67
rect 385 65 387 67
rect 667 65 669 67
rect 679 65 681 67
<< pdifct0 >>
rect 9 129 11 131
rect 40 136 42 138
rect 57 126 59 128
rect 74 136 76 138
rect 84 114 86 116
rect 105 136 107 138
rect 117 117 119 119
rect 140 136 142 138
rect 140 129 142 131
rect 152 128 154 130
rect 152 121 154 123
rect 162 136 164 138
rect 162 129 164 131
rect 194 136 196 138
rect 206 117 208 119
rect 229 136 231 138
rect 229 129 231 131
rect 241 128 243 130
rect 241 121 243 123
rect 251 136 253 138
rect 251 129 253 131
rect 272 129 274 131
rect 291 136 293 138
rect 326 128 328 130
rect 343 122 345 124
rect 360 128 362 130
rect 408 136 410 138
rect 621 137 623 139
rect 408 129 410 131
rect 427 129 429 131
rect 370 114 372 116
rect 444 123 446 125
rect 461 129 463 131
rect 491 129 493 131
rect 508 123 510 125
rect 525 129 527 131
rect 417 115 419 117
rect 555 129 557 131
rect 572 123 574 125
rect 589 129 591 131
rect 535 115 537 117
rect 639 130 641 132
rect 599 115 601 117
rect 660 115 662 117
rect 670 115 672 117
rect 680 119 682 121
rect 6 25 8 27
rect 16 29 18 31
rect 26 29 28 31
rect 87 29 89 31
rect 47 14 49 16
rect 151 29 153 31
rect 97 15 99 17
rect 114 21 116 23
rect 131 15 133 17
rect 269 29 271 31
rect 161 15 163 17
rect 178 21 180 23
rect 195 15 197 17
rect 225 15 227 17
rect 242 21 244 23
rect 316 30 318 32
rect 259 15 261 17
rect 278 15 280 17
rect 65 7 67 9
rect 278 8 280 10
rect 326 16 328 18
rect 343 22 345 24
rect 360 16 362 18
rect 395 8 397 10
rect 414 15 416 17
rect 435 15 437 17
rect 435 8 437 10
rect 445 23 447 25
rect 445 16 447 18
rect 457 15 459 17
rect 457 8 459 10
rect 480 27 482 29
rect 492 8 494 10
rect 524 15 526 17
rect 524 8 526 10
rect 534 23 536 25
rect 534 16 536 18
rect 546 15 548 17
rect 546 8 548 10
rect 569 27 571 29
rect 581 8 583 10
rect 602 30 604 32
rect 612 8 614 10
rect 629 18 631 20
rect 646 8 648 10
rect 677 15 679 17
<< pdifct1 >>
rect 30 129 32 131
rect 20 121 22 123
rect 20 114 22 116
rect 94 124 96 126
rect 94 117 96 119
rect 172 121 174 123
rect 172 114 174 116
rect 183 124 185 126
rect 183 117 185 119
rect 261 121 263 123
rect 261 114 263 116
rect 302 126 304 128
rect 302 119 304 121
rect 316 122 318 124
rect 389 130 391 132
rect 471 123 473 125
rect 481 123 483 125
rect 545 123 547 125
rect 609 128 611 130
rect 650 115 652 117
rect 36 29 38 31
rect 77 16 79 18
rect 141 21 143 23
rect 205 21 207 23
rect 215 21 217 23
rect 297 14 299 16
rect 370 22 372 24
rect 384 25 386 27
rect 384 18 386 20
rect 425 30 427 32
rect 425 23 427 25
rect 503 27 505 29
rect 503 20 505 22
rect 514 30 516 32
rect 514 23 516 25
rect 592 27 594 29
rect 592 20 594 22
rect 666 30 668 32
rect 666 23 668 25
rect 656 15 658 17
<< alu0 >>
rect 7 131 13 138
rect 38 136 40 138
rect 42 136 44 138
rect 38 135 44 136
rect 73 136 74 138
rect 76 136 77 138
rect 73 134 77 136
rect 103 136 105 138
rect 107 136 109 138
rect 103 135 109 136
rect 138 136 140 138
rect 142 136 144 138
rect 7 129 9 131
rect 11 129 13 131
rect 7 128 13 129
rect 48 128 61 129
rect 19 112 20 119
rect 5 95 9 97
rect 5 93 6 95
rect 8 93 9 95
rect 19 94 20 100
rect 5 82 9 93
rect 48 126 57 128
rect 59 126 61 128
rect 48 125 61 126
rect 36 121 52 125
rect 36 104 40 121
rect 138 131 144 136
rect 160 136 162 138
rect 164 136 166 138
rect 138 129 140 131
rect 142 129 144 131
rect 138 128 144 129
rect 151 130 155 132
rect 151 128 152 130
rect 154 128 155 130
rect 160 131 166 136
rect 192 136 194 138
rect 196 136 198 138
rect 192 135 198 136
rect 227 136 229 138
rect 231 136 233 138
rect 160 129 162 131
rect 164 129 166 131
rect 160 128 166 129
rect 227 131 233 136
rect 249 136 251 138
rect 253 136 255 138
rect 227 129 229 131
rect 231 129 233 131
rect 227 128 233 129
rect 240 130 244 132
rect 240 128 241 130
rect 243 128 244 130
rect 249 131 255 136
rect 289 136 291 138
rect 293 136 295 138
rect 289 135 295 136
rect 249 129 251 131
rect 253 129 255 131
rect 249 128 255 129
rect 270 131 287 132
rect 270 129 272 131
rect 274 129 287 131
rect 270 128 287 129
rect 108 124 132 128
rect 151 124 155 128
rect 60 117 64 119
rect 43 108 44 114
rect 60 115 61 117
rect 63 116 88 117
rect 63 115 84 116
rect 60 114 84 115
rect 86 114 88 116
rect 60 113 88 114
rect 35 102 40 104
rect 60 103 64 113
rect 35 100 36 102
rect 38 100 40 102
rect 53 101 64 103
rect 35 98 50 100
rect 36 96 50 98
rect 53 99 54 101
rect 56 99 64 101
rect 53 97 64 99
rect 39 90 43 92
rect 39 88 40 90
rect 42 88 43 90
rect 39 82 43 88
rect 46 91 50 96
rect 84 93 88 113
rect 72 92 78 93
rect 46 90 61 91
rect 46 88 57 90
rect 59 88 61 90
rect 46 87 61 88
rect 72 90 74 92
rect 76 90 78 92
rect 72 82 78 90
rect 82 92 88 93
rect 82 90 84 92
rect 86 90 88 92
rect 82 89 88 90
rect 106 120 112 124
rect 128 123 168 124
rect 128 121 152 123
rect 154 121 168 123
rect 106 110 110 120
rect 116 119 120 121
rect 128 120 168 121
rect 116 117 117 119
rect 119 117 120 119
rect 116 116 120 117
rect 106 108 107 110
rect 109 108 110 110
rect 106 106 110 108
rect 113 112 120 116
rect 113 101 117 112
rect 156 107 160 112
rect 156 105 157 107
rect 159 105 160 107
rect 99 100 117 101
rect 99 98 101 100
rect 103 99 117 100
rect 103 98 128 99
rect 99 97 124 98
rect 113 96 124 97
rect 126 96 128 98
rect 113 95 128 96
rect 133 98 137 100
rect 133 96 134 98
rect 136 96 137 98
rect 133 91 137 96
rect 112 90 134 91
rect 103 87 107 89
rect 112 88 114 90
rect 116 89 134 90
rect 136 89 137 91
rect 116 88 137 89
rect 112 87 137 88
rect 156 103 160 105
rect 164 109 168 120
rect 164 107 170 109
rect 164 105 167 107
rect 169 105 170 107
rect 164 103 170 105
rect 164 100 168 103
rect 148 96 168 100
rect 148 92 152 96
rect 144 91 152 92
rect 146 89 152 91
rect 144 88 152 89
rect 197 124 221 128
rect 240 124 244 128
rect 195 120 201 124
rect 217 123 257 124
rect 217 121 241 123
rect 243 121 257 123
rect 195 110 199 120
rect 205 119 209 121
rect 217 120 257 121
rect 205 117 206 119
rect 208 117 209 119
rect 205 116 209 117
rect 195 108 196 110
rect 198 108 199 110
rect 195 106 199 108
rect 202 112 209 116
rect 202 101 206 112
rect 245 107 249 112
rect 245 105 246 107
rect 248 105 249 107
rect 188 100 206 101
rect 188 98 190 100
rect 192 99 206 100
rect 192 98 217 99
rect 188 97 213 98
rect 202 96 213 97
rect 215 96 217 98
rect 202 95 217 96
rect 222 98 226 100
rect 222 96 223 98
rect 225 96 226 98
rect 222 91 226 96
rect 245 103 249 105
rect 253 109 257 120
rect 283 124 287 128
rect 283 120 298 124
rect 253 107 259 109
rect 253 105 256 107
rect 258 105 259 107
rect 253 103 259 105
rect 253 100 257 103
rect 237 96 257 100
rect 237 92 241 96
rect 273 111 279 112
rect 294 107 298 120
rect 301 117 302 128
rect 324 130 330 138
rect 324 128 326 130
rect 328 128 330 130
rect 324 127 330 128
rect 358 130 364 138
rect 407 136 408 138
rect 410 136 411 138
rect 358 128 360 130
rect 362 128 364 130
rect 358 127 364 128
rect 294 105 295 107
rect 297 105 298 107
rect 294 99 298 105
rect 280 98 298 99
rect 280 96 282 98
rect 284 96 298 98
rect 280 95 298 96
rect 341 124 347 125
rect 330 122 343 124
rect 345 122 347 124
rect 330 120 347 122
rect 407 131 411 136
rect 407 129 408 131
rect 410 129 411 131
rect 201 90 223 91
rect 192 87 196 89
rect 201 88 203 90
rect 205 89 223 90
rect 225 89 226 91
rect 205 88 226 89
rect 231 91 241 92
rect 231 89 233 91
rect 235 89 241 91
rect 231 88 241 89
rect 330 117 334 120
rect 321 113 334 117
rect 346 116 374 117
rect 321 99 325 113
rect 346 115 370 116
rect 346 113 347 115
rect 349 114 370 115
rect 372 114 374 116
rect 349 113 374 114
rect 346 101 350 113
rect 339 99 350 101
rect 321 97 322 99
rect 324 97 336 99
rect 321 95 336 97
rect 339 97 340 99
rect 342 97 350 99
rect 339 95 350 97
rect 201 87 226 88
rect 325 90 329 92
rect 325 88 326 90
rect 328 88 329 90
rect 103 85 104 87
rect 106 85 107 87
rect 192 85 193 87
rect 195 85 196 87
rect 270 85 276 86
rect 103 82 107 85
rect 159 84 165 85
rect 159 82 161 84
rect 163 82 165 84
rect 192 82 196 85
rect 248 84 254 85
rect 248 82 250 84
rect 252 82 254 84
rect 270 83 272 85
rect 274 83 276 85
rect 270 82 276 83
rect 289 85 295 86
rect 289 83 291 85
rect 293 83 295 85
rect 289 82 295 83
rect 325 82 329 88
rect 332 91 336 95
rect 370 91 374 113
rect 407 127 411 129
rect 425 131 431 139
rect 425 129 427 131
rect 429 129 431 131
rect 425 128 431 129
rect 459 131 465 139
rect 459 129 461 131
rect 463 129 465 131
rect 459 128 465 129
rect 489 131 495 139
rect 489 129 491 131
rect 493 129 495 131
rect 489 128 495 129
rect 523 131 529 139
rect 523 129 525 131
rect 527 129 529 131
rect 523 128 529 129
rect 553 131 559 139
rect 553 129 555 131
rect 557 129 559 131
rect 553 128 559 129
rect 587 131 593 139
rect 619 137 621 139
rect 623 137 625 139
rect 619 136 625 137
rect 587 129 589 131
rect 591 129 593 131
rect 587 128 593 129
rect 442 125 448 126
rect 442 123 444 125
rect 446 123 459 125
rect 442 121 459 123
rect 455 118 459 121
rect 415 117 443 118
rect 415 115 417 117
rect 419 116 443 117
rect 419 115 440 116
rect 415 114 440 115
rect 442 114 443 116
rect 332 90 347 91
rect 332 88 343 90
rect 345 88 347 90
rect 332 87 347 88
rect 358 90 364 91
rect 358 88 360 90
rect 362 88 364 90
rect 358 82 364 88
rect 368 90 374 91
rect 368 88 370 90
rect 372 88 374 90
rect 368 87 374 88
rect 385 97 389 99
rect 385 95 386 97
rect 388 95 389 97
rect 385 83 389 95
rect 406 97 411 99
rect 406 95 407 97
rect 409 95 411 97
rect 406 93 411 95
rect 407 83 411 93
rect 415 92 419 114
rect 439 102 443 114
rect 455 114 468 118
rect 439 100 450 102
rect 464 100 468 114
rect 439 98 447 100
rect 449 98 450 100
rect 439 96 450 98
rect 453 98 465 100
rect 467 98 468 100
rect 453 96 468 98
rect 453 92 457 96
rect 415 91 421 92
rect 415 89 417 91
rect 419 89 421 91
rect 415 88 421 89
rect 425 91 431 92
rect 425 89 427 91
rect 429 89 431 91
rect 425 83 431 89
rect 442 91 457 92
rect 442 89 444 91
rect 446 89 457 91
rect 442 88 457 89
rect 460 91 464 93
rect 460 89 461 91
rect 463 89 464 91
rect 460 83 464 89
rect 506 125 512 126
rect 495 123 508 125
rect 510 123 512 125
rect 495 121 512 123
rect 570 125 576 126
rect 559 123 572 125
rect 574 123 576 125
rect 559 121 576 123
rect 623 132 643 133
rect 623 130 639 132
rect 641 130 643 132
rect 623 129 643 130
rect 495 118 499 121
rect 486 114 499 118
rect 511 117 539 118
rect 486 100 490 114
rect 511 116 535 117
rect 511 114 512 116
rect 514 115 535 116
rect 537 115 539 117
rect 514 114 539 115
rect 511 102 515 114
rect 504 100 515 102
rect 486 98 487 100
rect 489 98 501 100
rect 486 96 501 98
rect 504 98 505 100
rect 507 98 515 100
rect 504 96 515 98
rect 490 91 494 93
rect 490 89 491 91
rect 493 89 494 91
rect 490 83 494 89
rect 497 92 501 96
rect 535 92 539 114
rect 497 91 512 92
rect 497 89 508 91
rect 510 89 512 91
rect 497 88 512 89
rect 523 91 529 92
rect 523 89 525 91
rect 527 89 529 91
rect 523 83 529 89
rect 533 91 539 92
rect 533 89 535 91
rect 537 89 539 91
rect 533 88 539 89
rect 559 118 563 121
rect 550 114 563 118
rect 575 117 603 118
rect 550 100 554 114
rect 575 116 599 117
rect 575 114 576 116
rect 578 115 599 116
rect 601 115 603 117
rect 578 114 603 115
rect 575 102 579 114
rect 568 100 579 102
rect 550 98 551 100
rect 553 98 565 100
rect 550 96 565 98
rect 568 98 569 100
rect 571 98 579 100
rect 568 96 579 98
rect 554 91 558 93
rect 554 89 555 91
rect 557 89 558 91
rect 554 83 558 89
rect 561 92 565 96
rect 599 92 603 114
rect 561 91 576 92
rect 561 89 572 91
rect 574 89 576 91
rect 561 88 576 89
rect 587 91 593 92
rect 587 89 589 91
rect 591 89 593 91
rect 587 83 593 89
rect 597 91 603 92
rect 597 89 599 91
rect 601 89 603 91
rect 597 88 603 89
rect 611 126 612 129
rect 623 125 627 129
rect 615 121 627 125
rect 615 109 619 121
rect 615 107 616 109
rect 618 107 619 109
rect 615 102 619 107
rect 615 98 632 102
rect 617 94 623 95
rect 617 92 619 94
rect 621 92 623 94
rect 617 83 623 92
rect 628 94 632 98
rect 652 113 653 119
rect 656 118 660 139
rect 679 121 683 139
rect 679 119 680 121
rect 682 119 683 121
rect 656 117 664 118
rect 656 115 660 117
rect 662 115 664 117
rect 656 114 664 115
rect 668 117 674 118
rect 679 117 683 119
rect 668 115 670 117
rect 672 115 674 117
rect 668 109 674 115
rect 655 108 674 109
rect 655 106 657 108
rect 659 106 674 108
rect 655 105 674 106
rect 628 92 629 94
rect 631 92 632 94
rect 628 90 632 92
rect 637 94 643 95
rect 637 92 639 94
rect 641 92 643 94
rect 637 83 643 92
rect 652 94 653 96
rect 664 92 668 105
rect 664 91 683 92
rect 664 89 679 91
rect 681 89 683 91
rect 664 88 683 89
rect 5 57 24 58
rect 5 55 7 57
rect 9 55 24 57
rect 5 54 24 55
rect 20 41 24 54
rect 35 50 36 52
rect 45 54 51 63
rect 45 52 47 54
rect 49 52 51 54
rect 45 51 51 52
rect 56 54 60 56
rect 56 52 57 54
rect 59 52 60 54
rect 14 40 33 41
rect 14 38 29 40
rect 31 38 33 40
rect 14 37 33 38
rect 14 31 20 37
rect 14 29 16 31
rect 18 29 20 31
rect 5 27 9 29
rect 14 28 20 29
rect 24 31 32 32
rect 24 29 26 31
rect 28 29 32 31
rect 24 28 32 29
rect 5 25 6 27
rect 8 25 9 27
rect 5 7 9 25
rect 28 7 32 28
rect 35 27 36 33
rect 56 48 60 52
rect 65 54 71 63
rect 65 52 67 54
rect 69 52 71 54
rect 65 51 71 52
rect 56 44 73 48
rect 69 39 73 44
rect 69 37 70 39
rect 72 37 73 39
rect 69 25 73 37
rect 61 21 73 25
rect 61 17 65 21
rect 76 17 77 20
rect 85 57 91 58
rect 85 55 87 57
rect 89 55 91 57
rect 85 54 91 55
rect 95 57 101 63
rect 95 55 97 57
rect 99 55 101 57
rect 95 54 101 55
rect 112 57 127 58
rect 112 55 114 57
rect 116 55 127 57
rect 112 54 127 55
rect 85 32 89 54
rect 123 50 127 54
rect 130 57 134 63
rect 130 55 131 57
rect 133 55 134 57
rect 130 53 134 55
rect 109 48 120 50
rect 109 46 117 48
rect 119 46 120 48
rect 123 48 138 50
rect 123 46 135 48
rect 137 46 138 48
rect 109 44 120 46
rect 109 32 113 44
rect 85 31 110 32
rect 85 29 87 31
rect 89 30 110 31
rect 112 30 113 32
rect 89 29 113 30
rect 134 32 138 46
rect 85 28 113 29
rect 125 28 138 32
rect 125 25 129 28
rect 149 57 155 58
rect 149 55 151 57
rect 153 55 155 57
rect 149 54 155 55
rect 159 57 165 63
rect 159 55 161 57
rect 163 55 165 57
rect 159 54 165 55
rect 176 57 191 58
rect 176 55 178 57
rect 180 55 191 57
rect 176 54 191 55
rect 149 32 153 54
rect 187 50 191 54
rect 194 57 198 63
rect 194 55 195 57
rect 197 55 198 57
rect 194 53 198 55
rect 173 48 184 50
rect 173 46 181 48
rect 183 46 184 48
rect 187 48 202 50
rect 187 46 199 48
rect 201 46 202 48
rect 173 44 184 46
rect 173 32 177 44
rect 149 31 174 32
rect 149 29 151 31
rect 153 30 174 31
rect 176 30 177 32
rect 153 29 177 30
rect 198 32 202 46
rect 149 28 177 29
rect 189 28 202 32
rect 189 25 193 28
rect 45 16 65 17
rect 45 14 47 16
rect 49 14 65 16
rect 45 13 65 14
rect 112 23 129 25
rect 112 21 114 23
rect 116 21 129 23
rect 112 20 118 21
rect 176 23 193 25
rect 176 21 178 23
rect 180 21 193 23
rect 176 20 182 21
rect 224 57 228 63
rect 224 55 225 57
rect 227 55 228 57
rect 224 53 228 55
rect 231 57 246 58
rect 231 55 242 57
rect 244 55 246 57
rect 231 54 246 55
rect 257 57 263 63
rect 257 55 259 57
rect 261 55 263 57
rect 257 54 263 55
rect 267 57 273 58
rect 267 55 269 57
rect 271 55 273 57
rect 267 54 273 55
rect 231 50 235 54
rect 220 48 235 50
rect 220 46 221 48
rect 223 46 235 48
rect 238 48 249 50
rect 238 46 239 48
rect 241 46 249 48
rect 220 32 224 46
rect 238 44 249 46
rect 220 28 233 32
rect 245 32 249 44
rect 269 32 273 54
rect 277 53 281 63
rect 277 51 282 53
rect 277 49 279 51
rect 281 49 282 51
rect 277 47 282 49
rect 299 51 303 63
rect 299 49 300 51
rect 302 49 303 51
rect 299 47 303 49
rect 314 58 320 59
rect 314 56 316 58
rect 318 56 320 58
rect 314 55 320 56
rect 324 58 330 64
rect 324 56 326 58
rect 328 56 330 58
rect 324 55 330 56
rect 341 58 356 59
rect 341 56 343 58
rect 345 56 356 58
rect 341 55 356 56
rect 245 30 246 32
rect 248 31 273 32
rect 248 30 269 31
rect 245 29 269 30
rect 271 29 273 31
rect 245 28 273 29
rect 229 25 233 28
rect 229 23 246 25
rect 229 21 242 23
rect 244 21 246 23
rect 240 20 246 21
rect 95 17 101 18
rect 95 15 97 17
rect 99 15 101 17
rect 63 9 69 10
rect 63 7 65 9
rect 67 7 69 9
rect 95 7 101 15
rect 129 17 135 18
rect 129 15 131 17
rect 133 15 135 17
rect 129 7 135 15
rect 159 17 165 18
rect 159 15 161 17
rect 163 15 165 17
rect 159 7 165 15
rect 193 17 199 18
rect 193 15 195 17
rect 197 15 199 17
rect 193 7 199 15
rect 223 17 229 18
rect 223 15 225 17
rect 227 15 229 17
rect 223 7 229 15
rect 257 17 263 18
rect 257 15 259 17
rect 261 15 263 17
rect 257 7 263 15
rect 277 17 281 19
rect 314 33 318 55
rect 352 51 356 55
rect 359 58 363 64
rect 393 63 399 64
rect 393 61 395 63
rect 397 61 399 63
rect 393 60 399 61
rect 412 63 418 64
rect 412 61 414 63
rect 416 61 418 63
rect 434 62 436 64
rect 438 62 440 64
rect 434 61 440 62
rect 492 61 496 64
rect 523 62 525 64
rect 527 62 529 64
rect 523 61 529 62
rect 581 61 585 64
rect 412 60 418 61
rect 492 59 493 61
rect 495 59 496 61
rect 581 59 582 61
rect 584 59 585 61
rect 359 56 360 58
rect 362 56 363 58
rect 359 54 363 56
rect 462 58 487 59
rect 447 57 457 58
rect 447 55 453 57
rect 455 55 457 57
rect 447 54 457 55
rect 462 57 483 58
rect 462 55 463 57
rect 465 56 483 57
rect 485 56 487 58
rect 492 57 496 59
rect 465 55 487 56
rect 338 49 349 51
rect 338 47 346 49
rect 348 47 349 49
rect 352 49 367 51
rect 352 47 364 49
rect 366 47 367 49
rect 338 45 349 47
rect 338 33 342 45
rect 314 32 339 33
rect 314 30 316 32
rect 318 31 339 32
rect 341 31 342 33
rect 318 30 342 31
rect 363 33 367 47
rect 314 29 342 30
rect 354 29 367 33
rect 354 26 358 29
rect 277 15 278 17
rect 280 15 281 17
rect 277 10 281 15
rect 341 24 358 26
rect 341 22 343 24
rect 345 22 358 24
rect 341 21 347 22
rect 390 50 408 51
rect 390 48 404 50
rect 406 48 408 50
rect 390 47 408 48
rect 390 41 394 47
rect 390 39 391 41
rect 393 39 394 41
rect 324 18 330 19
rect 324 16 326 18
rect 328 16 330 18
rect 277 8 278 10
rect 280 8 281 10
rect 324 8 330 16
rect 358 18 364 19
rect 358 16 360 18
rect 362 16 364 18
rect 358 8 364 16
rect 386 18 387 29
rect 390 26 394 39
rect 409 34 415 35
rect 447 50 451 54
rect 431 46 451 50
rect 431 43 435 46
rect 429 41 435 43
rect 429 39 430 41
rect 432 39 435 41
rect 429 37 435 39
rect 390 22 405 26
rect 401 18 405 22
rect 431 26 435 37
rect 439 41 443 43
rect 462 50 466 55
rect 462 48 463 50
rect 465 48 466 50
rect 462 46 466 48
rect 471 50 486 51
rect 471 48 473 50
rect 475 49 486 50
rect 475 48 500 49
rect 471 47 496 48
rect 482 46 496 47
rect 498 46 500 48
rect 482 45 500 46
rect 439 39 440 41
rect 442 39 443 41
rect 439 34 443 39
rect 482 34 486 45
rect 479 30 486 34
rect 489 38 493 40
rect 489 36 490 38
rect 492 36 493 38
rect 479 29 483 30
rect 479 27 480 29
rect 482 27 483 29
rect 431 25 471 26
rect 479 25 483 27
rect 489 26 493 36
rect 431 23 445 25
rect 447 23 471 25
rect 431 22 471 23
rect 487 22 493 26
rect 444 18 448 22
rect 467 18 491 22
rect 536 57 544 58
rect 536 55 542 57
rect 536 54 544 55
rect 536 50 540 54
rect 520 46 540 50
rect 520 43 524 46
rect 518 41 524 43
rect 518 39 519 41
rect 521 39 524 41
rect 518 37 524 39
rect 520 26 524 37
rect 528 41 532 43
rect 551 58 576 59
rect 551 57 572 58
rect 551 55 552 57
rect 554 56 572 57
rect 574 56 576 58
rect 581 57 585 59
rect 554 55 576 56
rect 551 50 555 55
rect 551 48 552 50
rect 554 48 555 50
rect 551 46 555 48
rect 560 50 575 51
rect 560 48 562 50
rect 564 49 575 50
rect 564 48 589 49
rect 560 47 585 48
rect 571 46 585 47
rect 587 46 589 48
rect 571 45 589 46
rect 528 39 529 41
rect 531 39 532 41
rect 528 34 532 39
rect 571 34 575 45
rect 568 30 575 34
rect 578 38 582 40
rect 578 36 579 38
rect 581 36 582 38
rect 568 29 572 30
rect 568 27 569 29
rect 571 27 572 29
rect 520 25 560 26
rect 568 25 572 27
rect 578 26 582 36
rect 520 23 534 25
rect 536 23 560 25
rect 520 22 560 23
rect 576 22 582 26
rect 600 56 606 57
rect 600 54 602 56
rect 604 54 606 56
rect 600 53 606 54
rect 610 56 616 64
rect 610 54 612 56
rect 614 54 616 56
rect 627 58 642 59
rect 627 56 629 58
rect 631 56 642 58
rect 627 55 642 56
rect 610 53 616 54
rect 600 33 604 53
rect 638 50 642 55
rect 645 58 649 64
rect 645 56 646 58
rect 648 56 649 58
rect 645 54 649 56
rect 624 47 635 49
rect 624 45 632 47
rect 634 45 635 47
rect 638 48 652 50
rect 638 46 653 48
rect 624 43 635 45
rect 648 44 650 46
rect 652 44 653 46
rect 624 33 628 43
rect 648 42 653 44
rect 600 32 628 33
rect 600 30 602 32
rect 604 31 628 32
rect 604 30 625 31
rect 600 29 625 30
rect 627 29 628 31
rect 644 32 645 38
rect 624 27 628 29
rect 533 18 537 22
rect 556 18 580 22
rect 401 17 418 18
rect 401 15 414 17
rect 416 15 418 17
rect 401 14 418 15
rect 433 17 439 18
rect 433 15 435 17
rect 437 15 439 17
rect 393 10 399 11
rect 393 8 395 10
rect 397 8 399 10
rect 433 10 439 15
rect 444 16 445 18
rect 447 16 448 18
rect 444 14 448 16
rect 455 17 461 18
rect 455 15 457 17
rect 459 15 461 17
rect 433 8 435 10
rect 437 8 439 10
rect 455 10 461 15
rect 522 17 528 18
rect 522 15 524 17
rect 526 15 528 17
rect 455 8 457 10
rect 459 8 461 10
rect 490 10 496 11
rect 490 8 492 10
rect 494 8 496 10
rect 522 10 528 15
rect 533 16 534 18
rect 536 16 537 18
rect 533 14 537 16
rect 544 17 550 18
rect 544 15 546 17
rect 548 15 550 17
rect 522 8 524 10
rect 526 8 528 10
rect 544 10 550 15
rect 648 25 652 42
rect 636 21 652 25
rect 627 20 640 21
rect 627 18 629 20
rect 631 18 640 20
rect 679 53 683 64
rect 668 46 669 52
rect 679 51 680 53
rect 682 51 683 53
rect 679 49 683 51
rect 668 27 669 34
rect 627 17 640 18
rect 675 17 681 18
rect 675 15 677 17
rect 679 15 681 17
rect 544 8 546 10
rect 548 8 550 10
rect 579 10 585 11
rect 579 8 581 10
rect 583 8 585 10
rect 611 10 615 12
rect 611 8 612 10
rect 614 8 615 10
rect 644 10 650 11
rect 644 8 646 10
rect 648 8 650 10
rect 675 8 681 15
<< via1 >>
rect 6 105 8 107
rect 21 100 23 102
rect 29 105 31 107
rect 81 121 83 123
rect 49 113 51 115
rect 69 97 71 99
rect 152 113 154 115
rect 93 93 95 95
rect 141 96 143 98
rect 174 96 176 98
rect 182 113 184 115
rect 214 105 216 107
rect 370 129 372 131
rect 303 107 305 109
rect 271 96 273 98
rect 339 107 341 109
rect 360 96 362 98
rect 416 129 418 131
rect 536 128 538 130
rect 600 129 602 131
rect 401 122 403 124
rect 385 110 387 112
rect 409 114 411 116
rect 429 98 431 100
rect 452 107 454 109
rect 472 107 474 109
rect 500 107 502 109
rect 524 98 526 100
rect 544 98 546 100
rect 569 110 571 112
rect 592 97 594 99
rect 608 110 610 112
rect 632 123 634 125
rect 640 106 642 108
rect 665 123 667 125
rect 681 106 683 108
rect 649 97 651 99
rect 37 47 39 49
rect 5 38 7 40
rect 21 21 23 23
rect 46 38 48 40
rect 54 21 56 23
rect 78 34 80 36
rect 94 47 96 49
rect 117 34 119 36
rect 142 46 144 48
rect 162 46 164 48
rect 186 37 188 39
rect 214 37 216 39
rect 234 37 236 39
rect 257 46 259 48
rect 277 30 279 32
rect 301 34 303 36
rect 285 22 287 24
rect 86 15 88 17
rect 150 16 152 18
rect 270 15 272 17
rect 375 56 377 58
rect 326 48 328 50
rect 347 37 349 39
rect 415 48 417 50
rect 383 37 385 39
rect 316 15 318 17
rect 472 39 474 41
rect 504 31 506 33
rect 512 48 514 50
rect 545 48 547 50
rect 593 51 595 53
rect 534 31 536 33
rect 617 47 619 49
rect 637 31 639 33
rect 602 23 604 25
rect 657 39 659 41
rect 665 44 667 46
rect 680 39 682 41
<< via2 >>
rect 84 122 86 124
rect 178 96 180 98
rect 141 89 143 91
rect 623 114 625 116
rect 63 30 65 32
rect 371 58 373 60
rect 545 51 547 53
rect 508 48 510 50
rect 601 14 603 16
<< via3 >>
rect 84 129 86 131
rect 141 92 143 94
rect 371 55 373 57
rect 545 12 547 14
<< labels >>
rlabel alu1 510 68 510 68 5 Vss
rlabel alu1 510 4 510 4 5 Vdd
rlabel alu1 344 4 344 4 2 vdd
rlabel alu1 344 68 344 68 2 vss
rlabel alu1 445 79 445 79 4 vss
rlabel alu1 445 143 445 143 4 vdd
rlabel alu1 509 79 509 79 6 vss
rlabel alu1 509 143 509 143 6 vdd
rlabel alu1 573 143 573 143 6 vdd
rlabel alu1 573 79 573 79 6 vss
rlabel alu1 666 143 666 143 6 vdd
rlabel alu1 625 79 625 79 6 vss
rlabel alu1 625 143 625 143 6 vdd
rlabel space 605 78 645 146 1 or
rlabel space 647 78 687 146 1 and
rlabel space 408 78 605 146 1 4x1_mux
rlabel alu1 666 79 666 79 6 vss
rlabel space 377 0 688 76 1 fafs
rlabel space 312 0 376 76 1 shift_mux
rlabel alu1 398 78 398 78 6 vss
rlabel alu1 398 142 398 142 6 vdd
rlabel ab 383 77 412 146 1 decoder
rlabel alu1 536 133 536 133 1 s1
rlabel alu2 475 130 475 130 1 s0
rlabel alu1 178 78 178 78 1 Vss
rlabel alu1 178 142 178 142 1 Vdd
rlabel alu1 344 142 344 142 6 vdd
rlabel alu1 344 78 344 78 6 vss
rlabel alu1 243 67 243 67 8 vss
rlabel alu1 243 3 243 3 8 vdd
rlabel alu1 179 67 179 67 2 vss
rlabel alu1 179 3 179 3 2 vdd
rlabel alu1 115 3 115 3 2 vdd
rlabel alu1 115 67 115 67 2 vss
rlabel alu1 22 3 22 3 2 vdd
rlabel alu1 63 67 63 67 2 vss
rlabel alu1 63 3 63 3 2 vdd
rlabel space 43 0 83 68 5 or
rlabel space 1 0 41 68 5 and
rlabel space 83 0 280 68 5 4x1_mux
rlabel alu1 22 67 22 67 2 vss
rlabel space 0 70 311 146 5 fafs
rlabel space 312 70 376 146 5 shift_mux
rlabel alu1 290 68 290 68 2 vss
rlabel alu1 290 4 290 4 2 vdd
rlabel ab 276 0 305 69 5 decoder
rlabel alu1 152 13 152 13 5 s1
rlabel alu2 213 16 213 16 5 s0
rlabel alu1 371 35 371 35 1 COUT0
rlabel alu2 458 49 458 49 1 A0
rlabel alu2 546 47 546 47 1 CIN0
rlabel alu1 594 35 594 35 1 SUM0
rlabel via1 638 32 638 32 1 B0
rlabel alu1 602 15 602 15 1 BINV
rlabel alu1 481 114 481 114 1 OUT0
rlabel alu1 207 44 207 44 1 OUT1
rlabel polyct0 62 116 62 116 1 B1
rlabel alu1 86 131 86 131 1 BINV
rlabel via1 142 98 142 98 1 CIN1
rlabel alu2 230 97 230 97 1 A1
rlabel alu2 316 110 316 110 1 COUT1
<< end >>
