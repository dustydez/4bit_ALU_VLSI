magic
tech scmos
timestamp 1760167772
<< ab >>
rect 5 5 223 77
<< nwell >>
rect 0 37 228 82
<< pwell >>
rect 0 0 228 37
<< poly >>
rect 14 71 16 75
rect 37 68 39 73
rect 44 68 46 73
rect 62 71 64 75
rect 72 71 74 75
rect 82 71 84 75
rect 103 71 105 75
rect 27 59 29 64
rect 14 33 16 46
rect 27 43 29 46
rect 126 68 128 73
rect 133 68 135 73
rect 151 71 153 75
rect 161 71 163 75
rect 171 71 173 75
rect 192 71 194 75
rect 199 71 201 75
rect 116 59 118 64
rect 20 41 29 43
rect 20 39 22 41
rect 24 39 26 41
rect 37 40 39 43
rect 44 40 46 43
rect 62 40 64 43
rect 72 40 74 43
rect 82 40 84 43
rect 20 37 26 39
rect 14 31 20 33
rect 14 29 16 31
rect 18 29 20 31
rect 14 27 20 29
rect 14 24 16 27
rect 24 24 26 37
rect 34 38 40 40
rect 34 36 36 38
rect 38 36 40 38
rect 34 34 40 36
rect 44 38 66 40
rect 44 36 55 38
rect 57 36 62 38
rect 64 36 66 38
rect 44 34 66 36
rect 70 38 76 40
rect 70 36 72 38
rect 74 36 76 38
rect 70 34 76 36
rect 80 38 86 40
rect 80 36 82 38
rect 84 36 86 38
rect 80 34 86 36
rect 34 31 36 34
rect 44 31 46 34
rect 64 31 66 34
rect 71 31 73 34
rect 14 7 16 11
rect 24 9 26 14
rect 34 12 36 17
rect 44 12 46 17
rect 82 25 84 34
rect 103 33 105 46
rect 116 43 118 46
rect 212 61 214 66
rect 192 47 194 50
rect 188 45 194 47
rect 188 43 190 45
rect 192 43 194 45
rect 109 41 118 43
rect 109 39 111 41
rect 113 39 115 41
rect 126 40 128 43
rect 133 40 135 43
rect 151 40 153 43
rect 161 40 163 43
rect 171 40 173 43
rect 188 41 194 43
rect 109 37 115 39
rect 103 31 109 33
rect 103 29 105 31
rect 107 29 109 31
rect 103 27 109 29
rect 103 24 105 27
rect 113 24 115 37
rect 123 38 129 40
rect 123 36 125 38
rect 127 36 129 38
rect 123 34 129 36
rect 133 38 155 40
rect 133 36 144 38
rect 146 36 151 38
rect 153 36 155 38
rect 133 34 155 36
rect 159 38 165 40
rect 159 36 161 38
rect 163 36 165 38
rect 159 34 165 36
rect 169 38 175 40
rect 169 36 171 38
rect 173 36 175 38
rect 169 34 175 36
rect 123 31 125 34
rect 133 31 135 34
rect 153 31 155 34
rect 160 31 162 34
rect 64 7 66 11
rect 71 7 73 11
rect 82 7 84 11
rect 103 7 105 11
rect 113 9 115 14
rect 123 12 125 17
rect 133 12 135 17
rect 171 25 173 34
rect 192 31 194 41
rect 199 40 201 50
rect 212 40 214 43
rect 198 38 204 40
rect 198 36 200 38
rect 202 36 204 38
rect 198 34 204 36
rect 208 38 214 40
rect 208 36 210 38
rect 212 36 214 38
rect 208 34 214 36
rect 202 31 204 34
rect 212 31 214 34
rect 192 20 194 25
rect 202 20 204 25
rect 212 17 214 22
rect 153 7 155 11
rect 160 7 162 11
rect 171 7 173 11
<< ndif >>
rect 29 24 34 31
rect 7 22 14 24
rect 7 20 9 22
rect 11 20 14 22
rect 7 18 14 20
rect 9 11 14 18
rect 16 18 24 24
rect 16 16 19 18
rect 21 16 24 18
rect 16 14 24 16
rect 26 21 34 24
rect 26 19 29 21
rect 31 19 34 21
rect 26 17 34 19
rect 36 29 44 31
rect 36 27 39 29
rect 41 27 44 29
rect 36 17 44 27
rect 46 29 53 31
rect 46 27 49 29
rect 51 27 53 29
rect 46 22 53 27
rect 59 24 64 31
rect 46 20 49 22
rect 51 20 53 22
rect 46 17 53 20
rect 57 22 64 24
rect 57 20 59 22
rect 61 20 64 22
rect 57 18 64 20
rect 26 14 31 17
rect 16 11 21 14
rect 59 11 64 18
rect 66 11 71 31
rect 73 25 80 31
rect 73 15 82 25
rect 73 13 76 15
rect 78 13 82 15
rect 73 11 82 13
rect 84 22 91 25
rect 118 24 123 31
rect 84 20 87 22
rect 89 20 91 22
rect 84 18 91 20
rect 96 22 103 24
rect 96 20 98 22
rect 100 20 103 22
rect 96 18 103 20
rect 84 11 89 18
rect 98 11 103 18
rect 105 18 113 24
rect 105 16 108 18
rect 110 16 113 18
rect 105 14 113 16
rect 115 21 123 24
rect 115 19 118 21
rect 120 19 123 21
rect 115 17 123 19
rect 125 29 133 31
rect 125 27 128 29
rect 130 27 133 29
rect 125 17 133 27
rect 135 29 142 31
rect 135 27 138 29
rect 140 27 142 29
rect 135 22 142 27
rect 148 24 153 31
rect 135 20 138 22
rect 140 20 142 22
rect 135 17 142 20
rect 146 22 153 24
rect 146 20 148 22
rect 150 20 153 22
rect 146 18 153 20
rect 115 14 120 17
rect 105 11 110 14
rect 148 11 153 18
rect 155 11 160 31
rect 162 25 169 31
rect 185 25 192 31
rect 194 29 202 31
rect 194 27 197 29
rect 199 27 202 29
rect 194 25 202 27
rect 204 25 212 31
rect 162 15 171 25
rect 162 13 165 15
rect 167 13 171 15
rect 162 11 171 13
rect 173 22 180 25
rect 173 20 176 22
rect 178 20 180 22
rect 173 18 180 20
rect 185 18 190 25
rect 206 22 212 25
rect 214 29 221 31
rect 214 27 217 29
rect 219 27 221 29
rect 214 25 221 27
rect 214 22 219 25
rect 206 18 210 22
rect 173 11 178 18
rect 185 16 191 18
rect 185 14 187 16
rect 189 14 191 16
rect 185 12 191 14
rect 204 16 210 18
rect 204 14 206 16
rect 208 14 210 16
rect 204 12 210 14
<< pdif >>
rect 9 59 14 71
rect 7 57 14 59
rect 7 55 9 57
rect 11 55 14 57
rect 7 50 14 55
rect 7 48 9 50
rect 11 48 14 50
rect 7 46 14 48
rect 16 69 25 71
rect 16 67 20 69
rect 22 67 25 69
rect 48 69 62 71
rect 48 68 55 69
rect 16 59 25 67
rect 32 59 37 68
rect 16 46 27 59
rect 29 50 37 59
rect 29 48 32 50
rect 34 48 37 50
rect 29 46 37 48
rect 32 43 37 46
rect 39 43 44 68
rect 46 67 55 68
rect 57 67 62 69
rect 46 62 62 67
rect 46 60 55 62
rect 57 60 62 62
rect 46 43 62 60
rect 64 61 72 71
rect 64 59 67 61
rect 69 59 72 61
rect 64 54 72 59
rect 64 52 67 54
rect 69 52 72 54
rect 64 43 72 52
rect 74 69 82 71
rect 74 67 77 69
rect 79 67 82 69
rect 74 62 82 67
rect 74 60 77 62
rect 79 60 82 62
rect 74 43 82 60
rect 84 56 89 71
rect 98 59 103 71
rect 96 57 103 59
rect 84 54 91 56
rect 84 52 87 54
rect 89 52 91 54
rect 84 47 91 52
rect 84 45 87 47
rect 89 45 91 47
rect 96 55 98 57
rect 100 55 103 57
rect 96 50 103 55
rect 96 48 98 50
rect 100 48 103 50
rect 96 46 103 48
rect 105 69 114 71
rect 105 67 109 69
rect 111 67 114 69
rect 137 69 151 71
rect 137 68 144 69
rect 105 59 114 67
rect 121 59 126 68
rect 105 46 116 59
rect 118 50 126 59
rect 118 48 121 50
rect 123 48 126 50
rect 118 46 126 48
rect 84 43 91 45
rect 121 43 126 46
rect 128 43 133 68
rect 135 67 144 68
rect 146 67 151 69
rect 135 62 151 67
rect 135 60 144 62
rect 146 60 151 62
rect 135 43 151 60
rect 153 61 161 71
rect 153 59 156 61
rect 158 59 161 61
rect 153 54 161 59
rect 153 52 156 54
rect 158 52 161 54
rect 153 43 161 52
rect 163 69 171 71
rect 163 67 166 69
rect 168 67 171 69
rect 163 62 171 67
rect 163 60 166 62
rect 168 60 171 62
rect 163 43 171 60
rect 173 56 178 71
rect 187 64 192 71
rect 185 62 192 64
rect 185 60 187 62
rect 189 60 192 62
rect 185 58 192 60
rect 173 54 180 56
rect 173 52 176 54
rect 178 52 180 54
rect 173 47 180 52
rect 187 50 192 58
rect 194 50 199 71
rect 201 69 210 71
rect 201 67 206 69
rect 208 67 210 69
rect 201 61 210 67
rect 201 50 212 61
rect 173 45 176 47
rect 178 45 180 47
rect 173 43 180 45
rect 204 43 212 50
rect 214 59 221 61
rect 214 57 217 59
rect 219 57 221 59
rect 214 52 221 57
rect 214 50 217 52
rect 219 50 221 52
rect 214 48 221 50
rect 214 43 219 48
<< alu1 >>
rect 3 72 225 77
rect 3 70 216 72
rect 218 70 225 72
rect 3 69 225 70
rect 7 59 20 63
rect 96 59 109 63
rect 217 63 221 64
rect 208 59 221 63
rect 7 57 12 59
rect 7 55 9 57
rect 11 55 12 57
rect 96 57 101 59
rect 7 50 12 55
rect 7 48 9 50
rect 11 48 12 50
rect 7 46 12 48
rect 7 43 11 46
rect 7 41 8 43
rect 10 41 11 43
rect 7 24 11 41
rect 38 43 76 47
rect 38 40 43 43
rect 35 38 43 40
rect 35 36 36 38
rect 38 36 43 38
rect 35 34 43 36
rect 53 38 68 39
rect 53 36 55 38
rect 57 36 62 38
rect 64 36 68 38
rect 53 35 68 36
rect 7 22 12 24
rect 55 26 59 35
rect 86 54 92 56
rect 86 52 87 54
rect 89 52 92 54
rect 86 47 92 52
rect 86 45 87 47
rect 89 45 92 47
rect 86 43 92 45
rect 88 30 92 43
rect 88 28 89 30
rect 91 28 92 30
rect 88 23 92 28
rect 7 20 9 22
rect 11 20 12 22
rect 7 18 12 20
rect 70 22 92 23
rect 70 20 87 22
rect 89 20 92 22
rect 70 19 92 20
rect 96 55 98 57
rect 100 55 101 57
rect 96 50 101 55
rect 96 48 98 50
rect 100 48 101 50
rect 96 46 101 48
rect 96 24 100 46
rect 127 43 165 47
rect 127 41 128 43
rect 130 41 132 43
rect 127 40 132 41
rect 124 38 132 40
rect 124 36 125 38
rect 127 36 132 38
rect 124 34 132 36
rect 142 38 157 39
rect 142 36 144 38
rect 146 36 151 38
rect 153 36 157 38
rect 142 35 157 36
rect 96 22 101 24
rect 144 26 148 35
rect 175 54 189 56
rect 175 52 176 54
rect 178 52 189 54
rect 175 47 181 52
rect 175 45 176 47
rect 178 45 181 47
rect 175 43 181 45
rect 185 47 189 52
rect 185 45 206 47
rect 185 43 190 45
rect 192 43 206 45
rect 177 23 181 43
rect 185 38 206 39
rect 185 36 200 38
rect 202 36 206 38
rect 185 35 206 36
rect 219 57 221 59
rect 217 52 221 57
rect 219 50 221 52
rect 185 30 189 35
rect 217 31 221 50
rect 185 28 186 30
rect 188 28 189 30
rect 185 26 189 28
rect 216 29 221 31
rect 216 27 217 29
rect 219 27 221 29
rect 216 25 221 27
rect 96 20 98 22
rect 100 20 101 22
rect 96 18 101 20
rect 159 22 181 23
rect 159 20 176 22
rect 178 20 181 22
rect 159 19 181 20
rect 3 12 225 13
rect 3 10 216 12
rect 218 10 225 12
rect 3 5 225 10
<< alu2 >>
rect 7 43 132 44
rect 7 41 8 43
rect 10 41 128 43
rect 130 41 132 43
rect 7 40 132 41
rect 88 30 189 31
rect 88 28 89 30
rect 91 28 186 30
rect 188 28 189 30
rect 88 27 189 28
<< ptie >>
rect 214 12 220 14
rect 214 10 216 12
rect 218 10 220 12
rect 214 8 220 10
<< ntie >>
rect 214 72 220 74
rect 214 70 216 72
rect 218 70 220 72
rect 214 68 220 70
<< nmos >>
rect 14 11 16 24
rect 24 14 26 24
rect 34 17 36 31
rect 44 17 46 31
rect 64 11 66 31
rect 71 11 73 31
rect 82 11 84 25
rect 103 11 105 24
rect 113 14 115 24
rect 123 17 125 31
rect 133 17 135 31
rect 153 11 155 31
rect 160 11 162 31
rect 192 25 194 31
rect 202 25 204 31
rect 171 11 173 25
rect 212 22 214 31
<< pmos >>
rect 14 46 16 71
rect 27 46 29 59
rect 37 43 39 68
rect 44 43 46 68
rect 62 43 64 71
rect 72 43 74 71
rect 82 43 84 71
rect 103 46 105 71
rect 116 46 118 59
rect 126 43 128 68
rect 133 43 135 68
rect 151 43 153 71
rect 161 43 163 71
rect 171 43 173 71
rect 192 50 194 71
rect 199 50 201 71
rect 212 43 214 61
<< polyct0 >>
rect 22 39 24 41
rect 16 29 18 31
rect 72 36 74 38
rect 82 36 84 38
rect 111 39 113 41
rect 105 29 107 31
rect 161 36 163 38
rect 171 36 173 38
rect 210 36 212 38
<< polyct1 >>
rect 36 36 38 38
rect 55 36 57 38
rect 62 36 64 38
rect 190 43 192 45
rect 125 36 127 38
rect 144 36 146 38
rect 151 36 153 38
rect 200 36 202 38
<< ndifct0 >>
rect 19 16 21 18
rect 29 19 31 21
rect 39 27 41 29
rect 49 27 51 29
rect 49 20 51 22
rect 59 20 61 22
rect 76 13 78 15
rect 108 16 110 18
rect 118 19 120 21
rect 128 27 130 29
rect 138 27 140 29
rect 138 20 140 22
rect 148 20 150 22
rect 197 27 199 29
rect 165 13 167 15
rect 187 14 189 16
rect 206 14 208 16
<< ndifct1 >>
rect 9 20 11 22
rect 87 20 89 22
rect 98 20 100 22
rect 176 20 178 22
rect 217 27 219 29
<< ntiect1 >>
rect 216 70 218 72
<< ptiect1 >>
rect 216 10 218 12
<< pdifct0 >>
rect 20 67 22 69
rect 32 48 34 50
rect 55 67 57 69
rect 55 60 57 62
rect 67 59 69 61
rect 67 52 69 54
rect 77 67 79 69
rect 77 60 79 62
rect 109 67 111 69
rect 121 48 123 50
rect 144 67 146 69
rect 144 60 146 62
rect 156 59 158 61
rect 156 52 158 54
rect 166 67 168 69
rect 166 60 168 62
rect 187 60 189 62
rect 206 67 208 69
<< pdifct1 >>
rect 9 55 11 57
rect 9 48 11 50
rect 87 52 89 54
rect 87 45 89 47
rect 98 55 100 57
rect 98 48 100 50
rect 176 52 178 54
rect 176 45 178 47
rect 217 57 219 59
rect 217 50 219 52
<< alu0 >>
rect 18 67 20 69
rect 22 67 24 69
rect 18 66 24 67
rect 53 67 55 69
rect 57 67 59 69
rect 53 62 59 67
rect 75 67 77 69
rect 79 67 81 69
rect 53 60 55 62
rect 57 60 59 62
rect 53 59 59 60
rect 66 61 70 63
rect 66 59 67 61
rect 69 59 70 61
rect 75 62 81 67
rect 107 67 109 69
rect 111 67 113 69
rect 107 66 113 67
rect 142 67 144 69
rect 146 67 148 69
rect 75 60 77 62
rect 79 60 81 62
rect 75 59 81 60
rect 142 62 148 67
rect 164 67 166 69
rect 168 67 170 69
rect 142 60 144 62
rect 146 60 148 62
rect 142 59 148 60
rect 155 61 159 63
rect 155 59 156 61
rect 158 59 159 61
rect 164 62 170 67
rect 204 67 206 69
rect 208 67 210 69
rect 204 66 210 67
rect 164 60 166 62
rect 168 60 170 62
rect 164 59 170 60
rect 185 62 202 63
rect 185 60 187 62
rect 189 60 202 62
rect 185 59 202 60
rect 23 55 47 59
rect 66 55 70 59
rect 21 51 27 55
rect 43 54 83 55
rect 43 52 67 54
rect 69 52 83 54
rect 21 41 25 51
rect 31 50 35 52
rect 43 51 83 52
rect 31 48 32 50
rect 34 48 35 50
rect 31 47 35 48
rect 21 39 22 41
rect 24 39 25 41
rect 21 37 25 39
rect 28 43 35 47
rect 28 32 32 43
rect 71 38 75 43
rect 71 36 72 38
rect 74 36 75 38
rect 14 31 32 32
rect 14 29 16 31
rect 18 30 32 31
rect 18 29 43 30
rect 14 28 39 29
rect 28 27 39 28
rect 41 27 43 29
rect 28 26 43 27
rect 48 29 52 31
rect 48 27 49 29
rect 51 27 52 29
rect 48 22 52 27
rect 71 34 75 36
rect 79 40 83 51
rect 79 38 85 40
rect 79 36 82 38
rect 84 36 85 38
rect 79 34 85 36
rect 79 31 83 34
rect 63 27 83 31
rect 63 23 67 27
rect 27 21 49 22
rect 18 18 22 20
rect 27 19 29 21
rect 31 20 49 21
rect 51 20 52 22
rect 31 19 52 20
rect 57 22 67 23
rect 57 20 59 22
rect 61 20 67 22
rect 57 19 67 20
rect 112 55 136 59
rect 155 55 159 59
rect 110 51 116 55
rect 132 54 172 55
rect 132 52 156 54
rect 158 52 172 54
rect 110 41 114 51
rect 120 50 124 52
rect 132 51 172 52
rect 120 48 121 50
rect 123 48 124 50
rect 120 47 124 48
rect 110 39 111 41
rect 113 39 114 41
rect 110 37 114 39
rect 117 43 124 47
rect 117 32 121 43
rect 160 38 164 43
rect 160 36 161 38
rect 163 36 164 38
rect 103 31 121 32
rect 103 29 105 31
rect 107 30 121 31
rect 107 29 132 30
rect 103 28 128 29
rect 117 27 128 28
rect 130 27 132 29
rect 117 26 132 27
rect 137 29 141 31
rect 137 27 138 29
rect 140 27 141 29
rect 137 22 141 27
rect 160 34 164 36
rect 168 40 172 51
rect 198 55 202 59
rect 198 51 213 55
rect 168 38 174 40
rect 168 36 171 38
rect 173 36 174 38
rect 168 34 174 36
rect 168 31 172 34
rect 152 27 172 31
rect 152 23 156 27
rect 188 42 194 43
rect 209 38 213 51
rect 216 48 217 59
rect 209 36 210 38
rect 212 36 213 38
rect 209 30 213 36
rect 195 29 213 30
rect 195 27 197 29
rect 199 27 213 29
rect 195 26 213 27
rect 116 21 138 22
rect 27 18 52 19
rect 107 18 111 20
rect 116 19 118 21
rect 120 20 138 21
rect 140 20 141 22
rect 120 19 141 20
rect 146 22 156 23
rect 146 20 148 22
rect 150 20 156 22
rect 146 19 156 20
rect 116 18 141 19
rect 18 16 19 18
rect 21 16 22 18
rect 107 16 108 18
rect 110 16 111 18
rect 185 16 191 17
rect 18 13 22 16
rect 74 15 80 16
rect 74 13 76 15
rect 78 13 80 15
rect 107 13 111 16
rect 163 15 169 16
rect 163 13 165 15
rect 167 13 169 15
rect 185 14 187 16
rect 189 14 191 16
rect 185 13 191 14
rect 204 16 210 17
rect 204 14 206 16
rect 208 14 210 16
rect 204 13 210 14
<< via1 >>
rect 8 41 10 43
rect 89 28 91 30
rect 128 41 130 43
rect 186 28 188 30
<< labels >>
rlabel alu2 55 44 55 44 1 B
rlabel alu1 59 37 59 37 1 A
rlabel alu1 149 37 149 37 1 Cin
rlabel alu1 99 60 99 60 1 Sum
rlabel alu1 219 44 219 44 1 Cout
rlabel alu1 118 73 118 73 1 Vdd
rlabel alu1 117 8 117 8 1 Vss
<< end >>
