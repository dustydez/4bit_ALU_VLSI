magic
tech scmos
timestamp 1761038610
<< ab >>
rect 157 221 266 293
rect 268 221 310 293
rect 312 221 375 293
rect 382 223 412 293
rect 413 292 490 293
rect 497 292 603 293
rect 609 292 686 293
rect 413 224 645 292
rect 646 224 686 292
rect 377 221 409 223
rect 279 217 311 219
rect 2 148 42 216
rect 43 148 275 216
rect 2 147 79 148
rect 85 147 191 148
rect 198 147 275 148
rect 276 147 306 217
rect 313 147 376 219
rect 378 147 420 219
rect 422 147 531 219
rect 157 74 266 146
rect 268 74 310 146
rect 312 74 375 146
rect 382 76 412 146
rect 413 145 490 146
rect 497 145 603 146
rect 609 145 686 146
rect 413 77 645 145
rect 646 77 686 145
rect 377 74 409 76
rect 279 70 311 72
rect 2 1 42 69
rect 43 1 275 69
rect 2 0 79 1
rect 85 0 191 1
rect 198 0 275 1
rect 276 0 306 70
rect 313 0 376 72
rect 378 0 420 72
rect 422 0 531 72
<< nwell >>
rect 0 254 688 293
rect 0 253 313 254
rect 352 253 380 254
rect 306 186 688 187
rect 0 107 688 186
rect 0 106 382 107
rect 308 39 336 40
rect 375 39 688 40
rect 0 0 688 39
<< pwell >>
rect 313 253 352 254
rect 380 253 688 254
rect 0 227 352 253
rect 372 227 688 253
rect 0 187 688 227
rect 0 186 306 187
rect 382 106 688 107
rect 0 66 688 106
rect 0 40 316 66
rect 336 40 688 66
rect 0 39 308 40
rect 336 39 375 40
<< poly >>
rect 35 287 37 291
rect 45 287 47 291
rect 52 287 54 291
rect 62 287 64 291
rect 69 287 71 291
rect 99 287 101 291
rect 15 277 17 282
rect 82 274 88 276
rect 82 272 84 274
rect 86 272 88 274
rect 15 256 17 259
rect 11 254 17 256
rect 11 252 13 254
rect 15 252 17 254
rect 11 250 17 252
rect 35 251 37 269
rect 45 261 47 271
rect 42 259 48 261
rect 42 257 44 259
rect 46 257 48 259
rect 42 255 48 257
rect 52 256 54 271
rect 62 266 64 271
rect 59 264 65 266
rect 59 262 61 264
rect 63 262 65 264
rect 59 260 65 262
rect 69 256 71 271
rect 79 270 88 272
rect 79 267 81 270
rect 122 284 124 289
rect 129 284 131 289
rect 147 287 149 291
rect 157 287 159 291
rect 167 287 169 291
rect 188 287 190 291
rect 112 275 114 280
rect 15 247 17 250
rect 34 249 40 251
rect 34 247 36 249
rect 38 247 40 249
rect 34 245 40 247
rect 35 242 37 245
rect 15 233 17 238
rect 45 241 47 255
rect 52 254 64 256
rect 52 248 58 250
rect 52 246 54 248
rect 56 246 58 248
rect 52 244 58 246
rect 52 241 54 244
rect 62 241 64 254
rect 69 254 75 256
rect 69 252 71 254
rect 73 252 75 254
rect 69 250 75 252
rect 69 241 71 250
rect 79 241 81 259
rect 99 249 101 262
rect 112 259 114 262
rect 211 284 213 289
rect 218 284 220 289
rect 236 287 238 291
rect 246 287 248 291
rect 256 287 258 291
rect 277 287 279 291
rect 284 287 286 291
rect 201 275 203 280
rect 105 257 114 259
rect 105 255 107 257
rect 109 255 111 257
rect 122 256 124 259
rect 129 256 131 259
rect 147 256 149 259
rect 157 256 159 259
rect 167 256 169 259
rect 105 253 111 255
rect 99 247 105 249
rect 99 245 101 247
rect 103 245 105 247
rect 99 243 105 245
rect 99 240 101 243
rect 109 240 111 253
rect 119 254 125 256
rect 119 252 121 254
rect 123 252 125 254
rect 119 250 125 252
rect 129 254 151 256
rect 129 252 140 254
rect 142 252 147 254
rect 149 252 151 254
rect 129 250 151 252
rect 155 254 161 256
rect 155 252 157 254
rect 159 252 161 254
rect 155 250 161 252
rect 165 254 171 256
rect 165 252 167 254
rect 169 252 171 254
rect 165 250 171 252
rect 119 247 121 250
rect 129 247 131 250
rect 149 247 151 250
rect 156 247 158 250
rect 35 228 37 233
rect 45 228 47 233
rect 52 228 54 233
rect 62 225 64 233
rect 69 229 71 233
rect 79 225 81 235
rect 62 223 81 225
rect 99 223 101 227
rect 109 225 111 230
rect 119 228 121 233
rect 129 228 131 233
rect 167 241 169 250
rect 188 249 190 262
rect 201 259 203 262
rect 394 287 396 291
rect 401 287 403 291
rect 297 277 299 282
rect 321 279 323 284
rect 331 279 333 284
rect 338 279 340 284
rect 348 279 350 284
rect 355 279 357 284
rect 277 263 279 266
rect 273 261 279 263
rect 273 259 275 261
rect 277 259 279 261
rect 194 257 203 259
rect 194 255 196 257
rect 198 255 200 257
rect 211 256 213 259
rect 218 256 220 259
rect 236 256 238 259
rect 246 256 248 259
rect 256 256 258 259
rect 273 257 279 259
rect 194 253 200 255
rect 188 247 194 249
rect 188 245 190 247
rect 192 245 194 247
rect 188 243 194 245
rect 188 240 190 243
rect 198 240 200 253
rect 208 254 214 256
rect 208 252 210 254
rect 212 252 214 254
rect 208 250 214 252
rect 218 254 240 256
rect 218 252 229 254
rect 231 252 236 254
rect 238 252 240 254
rect 218 250 240 252
rect 244 254 250 256
rect 244 252 246 254
rect 248 252 250 254
rect 244 250 250 252
rect 254 254 260 256
rect 254 252 256 254
rect 258 252 260 254
rect 254 250 260 252
rect 208 247 210 250
rect 218 247 220 250
rect 238 247 240 250
rect 245 247 247 250
rect 149 223 151 227
rect 156 223 158 227
rect 167 223 169 227
rect 188 223 190 227
rect 198 225 200 230
rect 208 228 210 233
rect 218 228 220 233
rect 256 241 258 250
rect 277 247 279 257
rect 284 256 286 266
rect 368 272 374 274
rect 368 270 370 272
rect 372 270 374 272
rect 297 256 299 259
rect 283 254 289 256
rect 283 252 285 254
rect 287 252 289 254
rect 283 250 289 252
rect 293 254 299 256
rect 293 252 295 254
rect 297 252 299 254
rect 293 250 299 252
rect 287 247 289 250
rect 297 247 299 250
rect 321 248 323 267
rect 331 258 333 267
rect 328 256 334 258
rect 328 254 330 256
rect 332 254 334 256
rect 328 252 334 254
rect 338 254 340 267
rect 348 264 350 267
rect 345 262 351 264
rect 345 260 347 262
rect 349 260 351 262
rect 345 258 351 260
rect 355 256 357 267
rect 365 268 374 270
rect 365 265 367 268
rect 627 288 629 292
rect 634 288 636 292
rect 432 280 434 285
rect 439 280 441 285
rect 449 280 451 285
rect 456 280 458 285
rect 466 280 468 285
rect 486 280 488 285
rect 496 280 498 285
rect 503 280 505 285
rect 513 280 515 285
rect 520 280 522 285
rect 550 280 552 285
rect 560 280 562 285
rect 567 280 569 285
rect 577 280 579 285
rect 584 280 586 285
rect 415 273 421 275
rect 415 271 417 273
rect 419 271 421 273
rect 415 269 424 271
rect 394 264 396 267
rect 391 262 397 264
rect 391 260 393 262
rect 395 260 397 262
rect 355 254 361 256
rect 338 252 350 254
rect 277 236 279 241
rect 287 236 289 241
rect 320 246 326 248
rect 320 244 322 246
rect 324 244 326 246
rect 320 242 326 244
rect 321 239 323 242
rect 331 239 333 252
rect 338 246 344 248
rect 338 244 340 246
rect 342 244 344 246
rect 338 242 344 244
rect 338 239 340 242
rect 348 239 350 252
rect 355 252 357 254
rect 359 252 361 254
rect 355 250 361 252
rect 355 239 357 250
rect 365 239 367 259
rect 391 258 397 260
rect 392 246 394 258
rect 401 255 403 267
rect 422 266 424 269
rect 533 273 539 275
rect 533 271 535 273
rect 537 271 539 273
rect 401 253 407 255
rect 401 251 403 253
rect 405 251 407 253
rect 401 249 407 251
rect 402 246 404 249
rect 422 240 424 260
rect 432 257 434 268
rect 439 265 441 268
rect 438 263 444 265
rect 438 261 440 263
rect 442 261 444 263
rect 438 259 444 261
rect 428 255 434 257
rect 449 255 451 268
rect 456 259 458 268
rect 428 253 430 255
rect 432 253 434 255
rect 428 251 434 253
rect 432 240 434 251
rect 439 253 451 255
rect 455 257 461 259
rect 455 255 457 257
rect 459 255 461 257
rect 455 253 461 255
rect 439 240 441 253
rect 445 247 451 249
rect 445 245 447 247
rect 449 245 451 247
rect 445 243 451 245
rect 449 240 451 243
rect 456 240 458 253
rect 466 249 468 268
rect 486 249 488 268
rect 496 259 498 268
rect 493 257 499 259
rect 493 255 495 257
rect 497 255 499 257
rect 493 253 499 255
rect 503 255 505 268
rect 513 265 515 268
rect 510 263 516 265
rect 510 261 512 263
rect 514 261 516 263
rect 510 259 516 261
rect 520 257 522 268
rect 530 269 539 271
rect 530 266 532 269
rect 614 279 616 283
rect 597 273 603 275
rect 597 271 599 273
rect 601 271 603 273
rect 520 255 526 257
rect 503 253 515 255
rect 463 247 469 249
rect 463 245 465 247
rect 467 245 469 247
rect 463 243 469 245
rect 485 247 491 249
rect 485 245 487 247
rect 489 245 491 247
rect 485 243 491 245
rect 466 240 468 243
rect 486 240 488 243
rect 496 240 498 253
rect 503 247 509 249
rect 503 245 505 247
rect 507 245 509 247
rect 503 243 509 245
rect 503 240 505 243
rect 513 240 515 253
rect 520 253 522 255
rect 524 253 526 255
rect 520 251 526 253
rect 520 240 522 251
rect 530 240 532 260
rect 550 249 552 268
rect 560 259 562 268
rect 557 257 563 259
rect 557 255 559 257
rect 561 255 563 257
rect 557 253 563 255
rect 567 255 569 268
rect 577 265 579 268
rect 574 263 580 265
rect 574 261 576 263
rect 578 261 580 263
rect 574 259 580 261
rect 584 257 586 268
rect 594 269 603 271
rect 594 266 596 269
rect 665 279 671 281
rect 665 277 667 279
rect 669 277 671 279
rect 655 272 657 277
rect 665 275 671 277
rect 584 255 590 257
rect 567 253 579 255
rect 549 247 555 249
rect 549 245 551 247
rect 553 245 555 247
rect 549 243 555 245
rect 550 240 552 243
rect 560 240 562 253
rect 567 247 573 249
rect 567 245 569 247
rect 571 245 573 247
rect 567 243 573 245
rect 567 240 569 243
rect 577 240 579 253
rect 584 253 586 255
rect 588 253 590 255
rect 584 251 590 253
rect 584 240 586 251
rect 594 240 596 260
rect 614 258 616 267
rect 627 265 629 270
rect 624 263 630 265
rect 624 261 626 263
rect 628 261 630 263
rect 624 259 630 261
rect 614 256 620 258
rect 614 254 616 256
rect 618 254 620 256
rect 614 252 620 254
rect 614 243 616 252
rect 624 243 626 259
rect 634 257 636 270
rect 665 270 667 275
rect 675 270 677 275
rect 655 257 657 260
rect 665 257 667 260
rect 634 255 640 257
rect 634 253 636 255
rect 638 253 640 255
rect 634 251 640 253
rect 655 255 661 257
rect 655 253 657 255
rect 659 253 661 255
rect 665 254 669 257
rect 655 251 661 253
rect 634 243 636 251
rect 655 243 657 251
rect 297 233 299 238
rect 392 235 394 240
rect 402 235 404 240
rect 667 240 669 254
rect 675 249 677 260
rect 674 247 680 249
rect 674 245 676 247
rect 678 245 680 247
rect 674 243 680 245
rect 674 240 676 243
rect 321 228 323 233
rect 331 228 333 233
rect 338 228 340 233
rect 238 223 240 227
rect 245 223 247 227
rect 256 223 258 227
rect 348 225 350 233
rect 355 229 357 233
rect 365 225 367 233
rect 348 223 367 225
rect 422 226 424 234
rect 432 230 434 234
rect 439 226 441 234
rect 449 229 451 234
rect 456 229 458 234
rect 466 229 468 234
rect 486 229 488 234
rect 496 229 498 234
rect 503 229 505 234
rect 422 224 441 226
rect 513 226 515 234
rect 520 230 522 234
rect 530 226 532 234
rect 550 229 552 234
rect 560 229 562 234
rect 567 229 569 234
rect 513 224 532 226
rect 577 226 579 234
rect 584 230 586 234
rect 594 226 596 234
rect 614 233 616 237
rect 624 233 626 237
rect 634 233 636 237
rect 655 233 657 237
rect 577 224 596 226
rect 667 226 669 231
rect 674 226 676 231
rect 12 209 14 214
rect 19 209 21 214
rect 92 214 111 216
rect 31 203 33 207
rect 52 203 54 207
rect 62 203 64 207
rect 72 203 74 207
rect 92 206 94 214
rect 102 206 104 210
rect 109 206 111 214
rect 156 214 175 216
rect 119 206 121 211
rect 126 206 128 211
rect 136 206 138 211
rect 156 206 158 214
rect 166 206 168 210
rect 173 206 175 214
rect 247 214 266 216
rect 183 206 185 211
rect 190 206 192 211
rect 200 206 202 211
rect 220 206 222 211
rect 230 206 232 211
rect 237 206 239 211
rect 247 206 249 214
rect 254 206 256 210
rect 264 206 266 214
rect 321 215 340 217
rect 321 207 323 215
rect 331 207 333 211
rect 338 207 340 215
rect 430 213 432 217
rect 441 213 443 217
rect 448 213 450 217
rect 348 207 350 212
rect 355 207 357 212
rect 365 207 367 212
rect 12 197 14 200
rect 8 195 14 197
rect 8 193 10 195
rect 12 193 14 195
rect 8 191 14 193
rect 11 180 13 191
rect 19 186 21 200
rect 284 200 286 205
rect 294 200 296 205
rect 389 202 391 207
rect 31 189 33 197
rect 52 189 54 197
rect 27 187 33 189
rect 19 183 23 186
rect 27 185 29 187
rect 31 185 33 187
rect 27 183 33 185
rect 48 187 54 189
rect 48 185 50 187
rect 52 185 54 187
rect 48 183 54 185
rect 21 180 23 183
rect 31 180 33 183
rect 11 165 13 170
rect 21 165 23 170
rect 52 170 54 183
rect 62 181 64 197
rect 72 188 74 197
rect 68 186 74 188
rect 68 184 70 186
rect 72 184 74 186
rect 68 182 74 184
rect 58 179 64 181
rect 58 177 60 179
rect 62 177 64 179
rect 58 175 64 177
rect 59 170 61 175
rect 72 173 74 182
rect 92 180 94 200
rect 102 189 104 200
rect 98 187 104 189
rect 98 185 100 187
rect 102 185 104 187
rect 109 187 111 200
rect 119 197 121 200
rect 115 195 121 197
rect 115 193 117 195
rect 119 193 121 195
rect 115 191 121 193
rect 126 187 128 200
rect 136 197 138 200
rect 133 195 139 197
rect 133 193 135 195
rect 137 193 139 195
rect 133 191 139 193
rect 109 185 121 187
rect 98 183 104 185
rect 17 163 23 165
rect 31 163 33 168
rect 17 161 19 163
rect 21 161 23 163
rect 17 159 23 161
rect 92 171 94 174
rect 85 169 94 171
rect 102 172 104 183
rect 108 179 114 181
rect 108 177 110 179
rect 112 177 114 179
rect 108 175 114 177
rect 109 172 111 175
rect 119 172 121 185
rect 125 185 131 187
rect 125 183 127 185
rect 129 183 131 185
rect 125 181 131 183
rect 126 172 128 181
rect 136 172 138 191
rect 156 180 158 200
rect 166 189 168 200
rect 162 187 168 189
rect 162 185 164 187
rect 166 185 168 187
rect 173 187 175 200
rect 183 197 185 200
rect 179 195 185 197
rect 179 193 181 195
rect 183 193 185 195
rect 179 191 185 193
rect 190 187 192 200
rect 200 197 202 200
rect 220 197 222 200
rect 197 195 203 197
rect 197 193 199 195
rect 201 193 203 195
rect 197 191 203 193
rect 219 195 225 197
rect 219 193 221 195
rect 223 193 225 195
rect 219 191 225 193
rect 173 185 185 187
rect 162 183 168 185
rect 85 167 87 169
rect 89 167 91 169
rect 85 165 91 167
rect 72 157 74 161
rect 156 171 158 174
rect 149 169 158 171
rect 166 172 168 183
rect 172 179 178 181
rect 172 177 174 179
rect 176 177 178 179
rect 172 175 178 177
rect 173 172 175 175
rect 183 172 185 185
rect 189 185 195 187
rect 189 183 191 185
rect 193 183 195 185
rect 189 181 195 183
rect 190 172 192 181
rect 200 172 202 191
rect 220 172 222 191
rect 230 187 232 200
rect 237 197 239 200
rect 237 195 243 197
rect 237 193 239 195
rect 241 193 243 195
rect 237 191 243 193
rect 247 187 249 200
rect 227 185 233 187
rect 227 183 229 185
rect 231 183 233 185
rect 227 181 233 183
rect 237 185 249 187
rect 254 189 256 200
rect 254 187 260 189
rect 254 185 256 187
rect 258 185 260 187
rect 230 172 232 181
rect 237 172 239 185
rect 254 183 260 185
rect 244 179 250 181
rect 244 177 246 179
rect 248 177 250 179
rect 244 175 250 177
rect 247 172 249 175
rect 254 172 256 183
rect 264 180 266 200
rect 284 191 286 194
rect 281 189 287 191
rect 281 187 283 189
rect 285 187 287 189
rect 281 185 287 187
rect 149 167 151 169
rect 153 167 155 169
rect 149 165 155 167
rect 264 171 266 174
rect 285 173 287 185
rect 294 182 296 194
rect 291 180 297 182
rect 321 181 323 201
rect 331 190 333 201
rect 327 188 333 190
rect 327 186 329 188
rect 331 186 333 188
rect 338 188 340 201
rect 348 198 350 201
rect 344 196 350 198
rect 344 194 346 196
rect 348 194 350 196
rect 344 192 350 194
rect 355 188 357 201
rect 365 198 367 201
rect 362 196 368 198
rect 362 194 364 196
rect 366 194 368 196
rect 362 192 368 194
rect 399 199 401 204
rect 409 199 411 204
rect 338 186 350 188
rect 327 184 333 186
rect 291 178 293 180
rect 295 178 297 180
rect 291 176 297 178
rect 292 173 294 176
rect 264 169 273 171
rect 267 167 269 169
rect 271 167 273 169
rect 267 165 273 167
rect 102 155 104 160
rect 109 155 111 160
rect 119 155 121 160
rect 126 155 128 160
rect 136 155 138 160
rect 166 155 168 160
rect 173 155 175 160
rect 183 155 185 160
rect 190 155 192 160
rect 200 155 202 160
rect 220 155 222 160
rect 230 155 232 160
rect 237 155 239 160
rect 247 155 249 160
rect 254 155 256 160
rect 52 148 54 152
rect 59 148 61 152
rect 321 172 323 175
rect 314 170 323 172
rect 331 173 333 184
rect 337 180 343 182
rect 337 178 339 180
rect 341 178 343 180
rect 337 176 343 178
rect 338 173 340 176
rect 348 173 350 186
rect 354 186 360 188
rect 354 184 356 186
rect 358 184 360 186
rect 354 182 360 184
rect 355 173 357 182
rect 365 173 367 192
rect 389 190 391 193
rect 399 190 401 193
rect 389 188 395 190
rect 389 186 391 188
rect 393 186 395 188
rect 389 184 395 186
rect 399 188 405 190
rect 399 186 401 188
rect 403 186 405 188
rect 399 184 405 186
rect 389 181 391 184
rect 314 168 316 170
rect 318 168 320 170
rect 314 166 320 168
rect 402 174 404 184
rect 409 183 411 193
rect 430 190 432 199
rect 468 207 470 212
rect 478 207 480 212
rect 488 210 490 215
rect 498 213 500 217
rect 519 213 521 217
rect 530 213 532 217
rect 537 213 539 217
rect 441 190 443 193
rect 448 190 450 193
rect 468 190 470 193
rect 478 190 480 193
rect 428 188 434 190
rect 428 186 430 188
rect 432 186 434 188
rect 428 184 434 186
rect 438 188 444 190
rect 438 186 440 188
rect 442 186 444 188
rect 438 184 444 186
rect 448 188 470 190
rect 448 186 450 188
rect 452 186 457 188
rect 459 186 470 188
rect 448 184 470 186
rect 474 188 480 190
rect 474 186 476 188
rect 478 186 480 188
rect 474 184 480 186
rect 488 187 490 200
rect 498 197 500 200
rect 494 195 500 197
rect 494 193 496 195
rect 498 193 500 195
rect 494 191 500 193
rect 488 185 494 187
rect 409 181 415 183
rect 430 181 432 184
rect 440 181 442 184
rect 450 181 452 184
rect 468 181 470 184
rect 475 181 477 184
rect 488 183 490 185
rect 492 183 494 185
rect 485 181 494 183
rect 409 179 411 181
rect 413 179 415 181
rect 409 177 415 179
rect 409 174 411 177
rect 331 156 333 161
rect 338 156 340 161
rect 348 156 350 161
rect 355 156 357 161
rect 365 156 367 161
rect 389 158 391 163
rect 285 149 287 153
rect 292 149 294 153
rect 485 178 487 181
rect 498 178 500 191
rect 519 190 521 199
rect 557 207 559 212
rect 567 207 569 212
rect 577 210 579 215
rect 587 213 589 217
rect 607 215 626 217
rect 607 205 609 215
rect 617 207 619 211
rect 624 207 626 215
rect 634 207 636 212
rect 641 207 643 212
rect 651 207 653 212
rect 530 190 532 193
rect 537 190 539 193
rect 557 190 559 193
rect 567 190 569 193
rect 517 188 523 190
rect 517 186 519 188
rect 521 186 523 188
rect 517 184 523 186
rect 527 188 533 190
rect 527 186 529 188
rect 531 186 533 188
rect 527 184 533 186
rect 537 188 559 190
rect 537 186 539 188
rect 541 186 546 188
rect 548 186 559 188
rect 537 184 559 186
rect 563 188 569 190
rect 563 186 565 188
rect 567 186 569 188
rect 563 184 569 186
rect 577 187 579 200
rect 587 197 589 200
rect 583 195 589 197
rect 583 193 585 195
rect 587 193 589 195
rect 583 191 589 193
rect 577 185 583 187
rect 519 181 521 184
rect 529 181 531 184
rect 539 181 541 184
rect 557 181 559 184
rect 564 181 566 184
rect 577 183 579 185
rect 581 183 583 185
rect 574 181 583 183
rect 485 160 487 165
rect 402 149 404 153
rect 409 149 411 153
rect 430 149 432 153
rect 440 149 442 153
rect 450 149 452 153
rect 468 151 470 156
rect 475 151 477 156
rect 574 178 576 181
rect 587 178 589 191
rect 607 181 609 199
rect 617 190 619 199
rect 613 188 619 190
rect 613 186 615 188
rect 617 186 619 188
rect 613 184 619 186
rect 624 186 626 199
rect 634 196 636 199
rect 630 194 636 196
rect 630 192 632 194
rect 634 192 636 194
rect 630 190 636 192
rect 624 184 636 186
rect 641 185 643 199
rect 671 202 673 207
rect 651 195 653 198
rect 648 193 654 195
rect 648 191 650 193
rect 652 191 654 193
rect 648 189 654 191
rect 671 190 673 193
rect 574 160 576 165
rect 498 149 500 153
rect 519 149 521 153
rect 529 149 531 153
rect 539 149 541 153
rect 557 151 559 156
rect 564 151 566 156
rect 607 170 609 173
rect 600 168 609 170
rect 617 169 619 184
rect 623 178 629 180
rect 623 176 625 178
rect 627 176 629 178
rect 623 174 629 176
rect 624 169 626 174
rect 634 169 636 184
rect 640 183 646 185
rect 640 181 642 183
rect 644 181 646 183
rect 640 179 646 181
rect 641 169 643 179
rect 651 171 653 189
rect 671 188 677 190
rect 671 186 673 188
rect 675 186 677 188
rect 671 184 677 186
rect 671 181 673 184
rect 600 166 602 168
rect 604 166 606 168
rect 600 164 606 166
rect 671 158 673 163
rect 587 149 589 153
rect 617 149 619 153
rect 624 149 626 153
rect 634 149 636 153
rect 641 149 643 153
rect 651 149 653 153
rect 35 140 37 144
rect 45 140 47 144
rect 52 140 54 144
rect 62 140 64 144
rect 69 140 71 144
rect 99 140 101 144
rect 15 130 17 135
rect 82 127 88 129
rect 82 125 84 127
rect 86 125 88 127
rect 15 109 17 112
rect 11 107 17 109
rect 11 105 13 107
rect 15 105 17 107
rect 11 103 17 105
rect 35 104 37 122
rect 45 114 47 124
rect 42 112 48 114
rect 42 110 44 112
rect 46 110 48 112
rect 42 108 48 110
rect 52 109 54 124
rect 62 119 64 124
rect 59 117 65 119
rect 59 115 61 117
rect 63 115 65 117
rect 59 113 65 115
rect 69 109 71 124
rect 79 123 88 125
rect 79 120 81 123
rect 122 137 124 142
rect 129 137 131 142
rect 147 140 149 144
rect 157 140 159 144
rect 167 140 169 144
rect 188 140 190 144
rect 112 128 114 133
rect 15 100 17 103
rect 34 102 40 104
rect 34 100 36 102
rect 38 100 40 102
rect 34 98 40 100
rect 35 95 37 98
rect 15 86 17 91
rect 45 94 47 108
rect 52 107 64 109
rect 52 101 58 103
rect 52 99 54 101
rect 56 99 58 101
rect 52 97 58 99
rect 52 94 54 97
rect 62 94 64 107
rect 69 107 75 109
rect 69 105 71 107
rect 73 105 75 107
rect 69 103 75 105
rect 69 94 71 103
rect 79 94 81 112
rect 99 102 101 115
rect 112 112 114 115
rect 211 137 213 142
rect 218 137 220 142
rect 236 140 238 144
rect 246 140 248 144
rect 256 140 258 144
rect 277 140 279 144
rect 284 140 286 144
rect 201 128 203 133
rect 105 110 114 112
rect 105 108 107 110
rect 109 108 111 110
rect 122 109 124 112
rect 129 109 131 112
rect 147 109 149 112
rect 157 109 159 112
rect 167 109 169 112
rect 105 106 111 108
rect 99 100 105 102
rect 99 98 101 100
rect 103 98 105 100
rect 99 96 105 98
rect 99 93 101 96
rect 109 93 111 106
rect 119 107 125 109
rect 119 105 121 107
rect 123 105 125 107
rect 119 103 125 105
rect 129 107 151 109
rect 129 105 140 107
rect 142 105 147 107
rect 149 105 151 107
rect 129 103 151 105
rect 155 107 161 109
rect 155 105 157 107
rect 159 105 161 107
rect 155 103 161 105
rect 165 107 171 109
rect 165 105 167 107
rect 169 105 171 107
rect 165 103 171 105
rect 119 100 121 103
rect 129 100 131 103
rect 149 100 151 103
rect 156 100 158 103
rect 35 81 37 86
rect 45 81 47 86
rect 52 81 54 86
rect 62 78 64 86
rect 69 82 71 86
rect 79 78 81 88
rect 62 76 81 78
rect 99 76 101 80
rect 109 78 111 83
rect 119 81 121 86
rect 129 81 131 86
rect 167 94 169 103
rect 188 102 190 115
rect 201 112 203 115
rect 394 140 396 144
rect 401 140 403 144
rect 297 130 299 135
rect 321 132 323 137
rect 331 132 333 137
rect 338 132 340 137
rect 348 132 350 137
rect 355 132 357 137
rect 277 116 279 119
rect 273 114 279 116
rect 273 112 275 114
rect 277 112 279 114
rect 194 110 203 112
rect 194 108 196 110
rect 198 108 200 110
rect 211 109 213 112
rect 218 109 220 112
rect 236 109 238 112
rect 246 109 248 112
rect 256 109 258 112
rect 273 110 279 112
rect 194 106 200 108
rect 188 100 194 102
rect 188 98 190 100
rect 192 98 194 100
rect 188 96 194 98
rect 188 93 190 96
rect 198 93 200 106
rect 208 107 214 109
rect 208 105 210 107
rect 212 105 214 107
rect 208 103 214 105
rect 218 107 240 109
rect 218 105 229 107
rect 231 105 236 107
rect 238 105 240 107
rect 218 103 240 105
rect 244 107 250 109
rect 244 105 246 107
rect 248 105 250 107
rect 244 103 250 105
rect 254 107 260 109
rect 254 105 256 107
rect 258 105 260 107
rect 254 103 260 105
rect 208 100 210 103
rect 218 100 220 103
rect 238 100 240 103
rect 245 100 247 103
rect 149 76 151 80
rect 156 76 158 80
rect 167 76 169 80
rect 188 76 190 80
rect 198 78 200 83
rect 208 81 210 86
rect 218 81 220 86
rect 256 94 258 103
rect 277 100 279 110
rect 284 109 286 119
rect 368 125 374 127
rect 368 123 370 125
rect 372 123 374 125
rect 297 109 299 112
rect 283 107 289 109
rect 283 105 285 107
rect 287 105 289 107
rect 283 103 289 105
rect 293 107 299 109
rect 293 105 295 107
rect 297 105 299 107
rect 293 103 299 105
rect 287 100 289 103
rect 297 100 299 103
rect 321 101 323 120
rect 331 111 333 120
rect 328 109 334 111
rect 328 107 330 109
rect 332 107 334 109
rect 328 105 334 107
rect 338 107 340 120
rect 348 117 350 120
rect 345 115 351 117
rect 345 113 347 115
rect 349 113 351 115
rect 345 111 351 113
rect 355 109 357 120
rect 365 121 374 123
rect 365 118 367 121
rect 627 141 629 145
rect 634 141 636 145
rect 432 133 434 138
rect 439 133 441 138
rect 449 133 451 138
rect 456 133 458 138
rect 466 133 468 138
rect 486 133 488 138
rect 496 133 498 138
rect 503 133 505 138
rect 513 133 515 138
rect 520 133 522 138
rect 550 133 552 138
rect 560 133 562 138
rect 567 133 569 138
rect 577 133 579 138
rect 584 133 586 138
rect 415 126 421 128
rect 415 124 417 126
rect 419 124 421 126
rect 415 122 424 124
rect 394 117 396 120
rect 391 115 397 117
rect 391 113 393 115
rect 395 113 397 115
rect 355 107 361 109
rect 338 105 350 107
rect 277 89 279 94
rect 287 89 289 94
rect 320 99 326 101
rect 320 97 322 99
rect 324 97 326 99
rect 320 95 326 97
rect 321 92 323 95
rect 331 92 333 105
rect 338 99 344 101
rect 338 97 340 99
rect 342 97 344 99
rect 338 95 344 97
rect 338 92 340 95
rect 348 92 350 105
rect 355 105 357 107
rect 359 105 361 107
rect 355 103 361 105
rect 355 92 357 103
rect 365 92 367 112
rect 391 111 397 113
rect 392 99 394 111
rect 401 108 403 120
rect 422 119 424 122
rect 533 126 539 128
rect 533 124 535 126
rect 537 124 539 126
rect 401 106 407 108
rect 401 104 403 106
rect 405 104 407 106
rect 401 102 407 104
rect 402 99 404 102
rect 422 93 424 113
rect 432 110 434 121
rect 439 118 441 121
rect 438 116 444 118
rect 438 114 440 116
rect 442 114 444 116
rect 438 112 444 114
rect 428 108 434 110
rect 449 108 451 121
rect 456 112 458 121
rect 428 106 430 108
rect 432 106 434 108
rect 428 104 434 106
rect 432 93 434 104
rect 439 106 451 108
rect 455 110 461 112
rect 455 108 457 110
rect 459 108 461 110
rect 455 106 461 108
rect 439 93 441 106
rect 445 100 451 102
rect 445 98 447 100
rect 449 98 451 100
rect 445 96 451 98
rect 449 93 451 96
rect 456 93 458 106
rect 466 102 468 121
rect 486 102 488 121
rect 496 112 498 121
rect 493 110 499 112
rect 493 108 495 110
rect 497 108 499 110
rect 493 106 499 108
rect 503 108 505 121
rect 513 118 515 121
rect 510 116 516 118
rect 510 114 512 116
rect 514 114 516 116
rect 510 112 516 114
rect 520 110 522 121
rect 530 122 539 124
rect 530 119 532 122
rect 614 132 616 136
rect 597 126 603 128
rect 597 124 599 126
rect 601 124 603 126
rect 520 108 526 110
rect 503 106 515 108
rect 463 100 469 102
rect 463 98 465 100
rect 467 98 469 100
rect 463 96 469 98
rect 485 100 491 102
rect 485 98 487 100
rect 489 98 491 100
rect 485 96 491 98
rect 466 93 468 96
rect 486 93 488 96
rect 496 93 498 106
rect 503 100 509 102
rect 503 98 505 100
rect 507 98 509 100
rect 503 96 509 98
rect 503 93 505 96
rect 513 93 515 106
rect 520 106 522 108
rect 524 106 526 108
rect 520 104 526 106
rect 520 93 522 104
rect 530 93 532 113
rect 550 102 552 121
rect 560 112 562 121
rect 557 110 563 112
rect 557 108 559 110
rect 561 108 563 110
rect 557 106 563 108
rect 567 108 569 121
rect 577 118 579 121
rect 574 116 580 118
rect 574 114 576 116
rect 578 114 580 116
rect 574 112 580 114
rect 584 110 586 121
rect 594 122 603 124
rect 594 119 596 122
rect 665 132 671 134
rect 665 130 667 132
rect 669 130 671 132
rect 655 125 657 130
rect 665 128 671 130
rect 584 108 590 110
rect 567 106 579 108
rect 549 100 555 102
rect 549 98 551 100
rect 553 98 555 100
rect 549 96 555 98
rect 550 93 552 96
rect 560 93 562 106
rect 567 100 573 102
rect 567 98 569 100
rect 571 98 573 100
rect 567 96 573 98
rect 567 93 569 96
rect 577 93 579 106
rect 584 106 586 108
rect 588 106 590 108
rect 584 104 590 106
rect 584 93 586 104
rect 594 93 596 113
rect 614 111 616 120
rect 627 118 629 123
rect 624 116 630 118
rect 624 114 626 116
rect 628 114 630 116
rect 624 112 630 114
rect 614 109 620 111
rect 614 107 616 109
rect 618 107 620 109
rect 614 105 620 107
rect 614 96 616 105
rect 624 96 626 112
rect 634 110 636 123
rect 665 123 667 128
rect 675 123 677 128
rect 655 110 657 113
rect 665 110 667 113
rect 634 108 640 110
rect 634 106 636 108
rect 638 106 640 108
rect 634 104 640 106
rect 655 108 661 110
rect 655 106 657 108
rect 659 106 661 108
rect 665 107 669 110
rect 655 104 661 106
rect 634 96 636 104
rect 655 96 657 104
rect 297 86 299 91
rect 392 88 394 93
rect 402 88 404 93
rect 667 93 669 107
rect 675 102 677 113
rect 674 100 680 102
rect 674 98 676 100
rect 678 98 680 100
rect 674 96 680 98
rect 674 93 676 96
rect 321 81 323 86
rect 331 81 333 86
rect 338 81 340 86
rect 238 76 240 80
rect 245 76 247 80
rect 256 76 258 80
rect 348 78 350 86
rect 355 82 357 86
rect 365 78 367 86
rect 348 76 367 78
rect 422 79 424 87
rect 432 83 434 87
rect 439 79 441 87
rect 449 82 451 87
rect 456 82 458 87
rect 466 82 468 87
rect 486 82 488 87
rect 496 82 498 87
rect 503 82 505 87
rect 422 77 441 79
rect 513 79 515 87
rect 520 83 522 87
rect 530 79 532 87
rect 550 82 552 87
rect 560 82 562 87
rect 567 82 569 87
rect 513 77 532 79
rect 577 79 579 87
rect 584 83 586 87
rect 594 79 596 87
rect 614 86 616 90
rect 624 86 626 90
rect 634 86 636 90
rect 655 86 657 90
rect 577 77 596 79
rect 667 79 669 84
rect 674 79 676 84
rect 12 62 14 67
rect 19 62 21 67
rect 92 67 111 69
rect 31 56 33 60
rect 52 56 54 60
rect 62 56 64 60
rect 72 56 74 60
rect 92 59 94 67
rect 102 59 104 63
rect 109 59 111 67
rect 156 67 175 69
rect 119 59 121 64
rect 126 59 128 64
rect 136 59 138 64
rect 156 59 158 67
rect 166 59 168 63
rect 173 59 175 67
rect 247 67 266 69
rect 183 59 185 64
rect 190 59 192 64
rect 200 59 202 64
rect 220 59 222 64
rect 230 59 232 64
rect 237 59 239 64
rect 247 59 249 67
rect 254 59 256 63
rect 264 59 266 67
rect 321 68 340 70
rect 321 60 323 68
rect 331 60 333 64
rect 338 60 340 68
rect 430 66 432 70
rect 441 66 443 70
rect 448 66 450 70
rect 348 60 350 65
rect 355 60 357 65
rect 365 60 367 65
rect 12 50 14 53
rect 8 48 14 50
rect 8 46 10 48
rect 12 46 14 48
rect 8 44 14 46
rect 11 33 13 44
rect 19 39 21 53
rect 284 53 286 58
rect 294 53 296 58
rect 389 55 391 60
rect 31 42 33 50
rect 52 42 54 50
rect 27 40 33 42
rect 19 36 23 39
rect 27 38 29 40
rect 31 38 33 40
rect 27 36 33 38
rect 48 40 54 42
rect 48 38 50 40
rect 52 38 54 40
rect 48 36 54 38
rect 21 33 23 36
rect 31 33 33 36
rect 11 18 13 23
rect 21 18 23 23
rect 52 23 54 36
rect 62 34 64 50
rect 72 41 74 50
rect 68 39 74 41
rect 68 37 70 39
rect 72 37 74 39
rect 68 35 74 37
rect 58 32 64 34
rect 58 30 60 32
rect 62 30 64 32
rect 58 28 64 30
rect 59 23 61 28
rect 72 26 74 35
rect 92 33 94 53
rect 102 42 104 53
rect 98 40 104 42
rect 98 38 100 40
rect 102 38 104 40
rect 109 40 111 53
rect 119 50 121 53
rect 115 48 121 50
rect 115 46 117 48
rect 119 46 121 48
rect 115 44 121 46
rect 126 40 128 53
rect 136 50 138 53
rect 133 48 139 50
rect 133 46 135 48
rect 137 46 139 48
rect 133 44 139 46
rect 109 38 121 40
rect 98 36 104 38
rect 17 16 23 18
rect 31 16 33 21
rect 17 14 19 16
rect 21 14 23 16
rect 17 12 23 14
rect 92 24 94 27
rect 85 22 94 24
rect 102 25 104 36
rect 108 32 114 34
rect 108 30 110 32
rect 112 30 114 32
rect 108 28 114 30
rect 109 25 111 28
rect 119 25 121 38
rect 125 38 131 40
rect 125 36 127 38
rect 129 36 131 38
rect 125 34 131 36
rect 126 25 128 34
rect 136 25 138 44
rect 156 33 158 53
rect 166 42 168 53
rect 162 40 168 42
rect 162 38 164 40
rect 166 38 168 40
rect 173 40 175 53
rect 183 50 185 53
rect 179 48 185 50
rect 179 46 181 48
rect 183 46 185 48
rect 179 44 185 46
rect 190 40 192 53
rect 200 50 202 53
rect 220 50 222 53
rect 197 48 203 50
rect 197 46 199 48
rect 201 46 203 48
rect 197 44 203 46
rect 219 48 225 50
rect 219 46 221 48
rect 223 46 225 48
rect 219 44 225 46
rect 173 38 185 40
rect 162 36 168 38
rect 85 20 87 22
rect 89 20 91 22
rect 85 18 91 20
rect 72 10 74 14
rect 156 24 158 27
rect 149 22 158 24
rect 166 25 168 36
rect 172 32 178 34
rect 172 30 174 32
rect 176 30 178 32
rect 172 28 178 30
rect 173 25 175 28
rect 183 25 185 38
rect 189 38 195 40
rect 189 36 191 38
rect 193 36 195 38
rect 189 34 195 36
rect 190 25 192 34
rect 200 25 202 44
rect 220 25 222 44
rect 230 40 232 53
rect 237 50 239 53
rect 237 48 243 50
rect 237 46 239 48
rect 241 46 243 48
rect 237 44 243 46
rect 247 40 249 53
rect 227 38 233 40
rect 227 36 229 38
rect 231 36 233 38
rect 227 34 233 36
rect 237 38 249 40
rect 254 42 256 53
rect 254 40 260 42
rect 254 38 256 40
rect 258 38 260 40
rect 230 25 232 34
rect 237 25 239 38
rect 254 36 260 38
rect 244 32 250 34
rect 244 30 246 32
rect 248 30 250 32
rect 244 28 250 30
rect 247 25 249 28
rect 254 25 256 36
rect 264 33 266 53
rect 284 44 286 47
rect 281 42 287 44
rect 281 40 283 42
rect 285 40 287 42
rect 281 38 287 40
rect 149 20 151 22
rect 153 20 155 22
rect 149 18 155 20
rect 264 24 266 27
rect 285 26 287 38
rect 294 35 296 47
rect 291 33 297 35
rect 321 34 323 54
rect 331 43 333 54
rect 327 41 333 43
rect 327 39 329 41
rect 331 39 333 41
rect 338 41 340 54
rect 348 51 350 54
rect 344 49 350 51
rect 344 47 346 49
rect 348 47 350 49
rect 344 45 350 47
rect 355 41 357 54
rect 365 51 367 54
rect 362 49 368 51
rect 362 47 364 49
rect 366 47 368 49
rect 362 45 368 47
rect 399 52 401 57
rect 409 52 411 57
rect 338 39 350 41
rect 327 37 333 39
rect 291 31 293 33
rect 295 31 297 33
rect 291 29 297 31
rect 292 26 294 29
rect 264 22 273 24
rect 267 20 269 22
rect 271 20 273 22
rect 267 18 273 20
rect 102 8 104 13
rect 109 8 111 13
rect 119 8 121 13
rect 126 8 128 13
rect 136 8 138 13
rect 166 8 168 13
rect 173 8 175 13
rect 183 8 185 13
rect 190 8 192 13
rect 200 8 202 13
rect 220 8 222 13
rect 230 8 232 13
rect 237 8 239 13
rect 247 8 249 13
rect 254 8 256 13
rect 52 1 54 5
rect 59 1 61 5
rect 321 25 323 28
rect 314 23 323 25
rect 331 26 333 37
rect 337 33 343 35
rect 337 31 339 33
rect 341 31 343 33
rect 337 29 343 31
rect 338 26 340 29
rect 348 26 350 39
rect 354 39 360 41
rect 354 37 356 39
rect 358 37 360 39
rect 354 35 360 37
rect 355 26 357 35
rect 365 26 367 45
rect 389 43 391 46
rect 399 43 401 46
rect 389 41 395 43
rect 389 39 391 41
rect 393 39 395 41
rect 389 37 395 39
rect 399 41 405 43
rect 399 39 401 41
rect 403 39 405 41
rect 399 37 405 39
rect 389 34 391 37
rect 314 21 316 23
rect 318 21 320 23
rect 314 19 320 21
rect 402 27 404 37
rect 409 36 411 46
rect 430 43 432 52
rect 468 60 470 65
rect 478 60 480 65
rect 488 63 490 68
rect 498 66 500 70
rect 519 66 521 70
rect 530 66 532 70
rect 537 66 539 70
rect 441 43 443 46
rect 448 43 450 46
rect 468 43 470 46
rect 478 43 480 46
rect 428 41 434 43
rect 428 39 430 41
rect 432 39 434 41
rect 428 37 434 39
rect 438 41 444 43
rect 438 39 440 41
rect 442 39 444 41
rect 438 37 444 39
rect 448 41 470 43
rect 448 39 450 41
rect 452 39 457 41
rect 459 39 470 41
rect 448 37 470 39
rect 474 41 480 43
rect 474 39 476 41
rect 478 39 480 41
rect 474 37 480 39
rect 488 40 490 53
rect 498 50 500 53
rect 494 48 500 50
rect 494 46 496 48
rect 498 46 500 48
rect 494 44 500 46
rect 488 38 494 40
rect 409 34 415 36
rect 430 34 432 37
rect 440 34 442 37
rect 450 34 452 37
rect 468 34 470 37
rect 475 34 477 37
rect 488 36 490 38
rect 492 36 494 38
rect 485 34 494 36
rect 409 32 411 34
rect 413 32 415 34
rect 409 30 415 32
rect 409 27 411 30
rect 331 9 333 14
rect 338 9 340 14
rect 348 9 350 14
rect 355 9 357 14
rect 365 9 367 14
rect 389 11 391 16
rect 285 2 287 6
rect 292 2 294 6
rect 485 31 487 34
rect 498 31 500 44
rect 519 43 521 52
rect 557 60 559 65
rect 567 60 569 65
rect 577 63 579 68
rect 587 66 589 70
rect 607 68 626 70
rect 607 58 609 68
rect 617 60 619 64
rect 624 60 626 68
rect 634 60 636 65
rect 641 60 643 65
rect 651 60 653 65
rect 530 43 532 46
rect 537 43 539 46
rect 557 43 559 46
rect 567 43 569 46
rect 517 41 523 43
rect 517 39 519 41
rect 521 39 523 41
rect 517 37 523 39
rect 527 41 533 43
rect 527 39 529 41
rect 531 39 533 41
rect 527 37 533 39
rect 537 41 559 43
rect 537 39 539 41
rect 541 39 546 41
rect 548 39 559 41
rect 537 37 559 39
rect 563 41 569 43
rect 563 39 565 41
rect 567 39 569 41
rect 563 37 569 39
rect 577 40 579 53
rect 587 50 589 53
rect 583 48 589 50
rect 583 46 585 48
rect 587 46 589 48
rect 583 44 589 46
rect 577 38 583 40
rect 519 34 521 37
rect 529 34 531 37
rect 539 34 541 37
rect 557 34 559 37
rect 564 34 566 37
rect 577 36 579 38
rect 581 36 583 38
rect 574 34 583 36
rect 485 13 487 18
rect 402 2 404 6
rect 409 2 411 6
rect 430 2 432 6
rect 440 2 442 6
rect 450 2 452 6
rect 468 4 470 9
rect 475 4 477 9
rect 574 31 576 34
rect 587 31 589 44
rect 607 34 609 52
rect 617 43 619 52
rect 613 41 619 43
rect 613 39 615 41
rect 617 39 619 41
rect 613 37 619 39
rect 624 39 626 52
rect 634 49 636 52
rect 630 47 636 49
rect 630 45 632 47
rect 634 45 636 47
rect 630 43 636 45
rect 624 37 636 39
rect 641 38 643 52
rect 671 55 673 60
rect 651 48 653 51
rect 648 46 654 48
rect 648 44 650 46
rect 652 44 654 46
rect 648 42 654 44
rect 671 43 673 46
rect 574 13 576 18
rect 498 2 500 6
rect 519 2 521 6
rect 529 2 531 6
rect 539 2 541 6
rect 557 4 559 9
rect 564 4 566 9
rect 607 23 609 26
rect 600 21 609 23
rect 617 22 619 37
rect 623 31 629 33
rect 623 29 625 31
rect 627 29 629 31
rect 623 27 629 29
rect 624 22 626 27
rect 634 22 636 37
rect 640 36 646 38
rect 640 34 642 36
rect 644 34 646 36
rect 640 32 646 34
rect 641 22 643 32
rect 651 24 653 42
rect 671 41 677 43
rect 671 39 673 41
rect 675 39 677 41
rect 671 37 677 39
rect 671 34 673 37
rect 600 19 602 21
rect 604 19 606 21
rect 600 17 606 19
rect 671 11 673 16
rect 587 2 589 6
rect 617 2 619 6
rect 624 2 626 6
rect 634 2 636 6
rect 641 2 643 6
rect 651 2 653 6
<< ndif >>
rect 4 242 15 247
rect 4 240 6 242
rect 8 240 15 242
rect 4 238 15 240
rect 17 245 24 247
rect 17 243 20 245
rect 22 243 24 245
rect 17 241 24 243
rect 17 238 22 241
rect 28 240 35 242
rect 28 238 30 240
rect 32 238 35 240
rect 28 236 35 238
rect 30 233 35 236
rect 37 241 42 242
rect 37 237 45 241
rect 37 235 40 237
rect 42 235 45 237
rect 37 233 45 235
rect 47 233 52 241
rect 54 237 62 241
rect 54 235 57 237
rect 59 235 62 237
rect 54 233 62 235
rect 64 233 69 241
rect 71 239 79 241
rect 71 237 74 239
rect 76 237 79 239
rect 71 235 79 237
rect 81 239 88 241
rect 114 240 119 247
rect 81 237 84 239
rect 86 237 88 239
rect 81 235 88 237
rect 92 238 99 240
rect 92 236 94 238
rect 96 236 99 238
rect 71 233 77 235
rect 92 234 99 236
rect 94 227 99 234
rect 101 234 109 240
rect 101 232 104 234
rect 106 232 109 234
rect 101 230 109 232
rect 111 237 119 240
rect 111 235 114 237
rect 116 235 119 237
rect 111 233 119 235
rect 121 245 129 247
rect 121 243 124 245
rect 126 243 129 245
rect 121 233 129 243
rect 131 245 138 247
rect 131 243 134 245
rect 136 243 138 245
rect 131 238 138 243
rect 144 240 149 247
rect 131 236 134 238
rect 136 236 138 238
rect 131 233 138 236
rect 142 238 149 240
rect 142 236 144 238
rect 146 236 149 238
rect 142 234 149 236
rect 111 230 116 233
rect 101 227 106 230
rect 144 227 149 234
rect 151 227 156 247
rect 158 241 165 247
rect 158 231 167 241
rect 158 229 161 231
rect 163 229 167 231
rect 158 227 167 229
rect 169 238 176 241
rect 203 240 208 247
rect 169 236 172 238
rect 174 236 176 238
rect 169 234 176 236
rect 181 238 188 240
rect 181 236 183 238
rect 185 236 188 238
rect 181 234 188 236
rect 169 227 174 234
rect 183 227 188 234
rect 190 234 198 240
rect 190 232 193 234
rect 195 232 198 234
rect 190 230 198 232
rect 200 237 208 240
rect 200 235 203 237
rect 205 235 208 237
rect 200 233 208 235
rect 210 245 218 247
rect 210 243 213 245
rect 215 243 218 245
rect 210 233 218 243
rect 220 245 227 247
rect 220 243 223 245
rect 225 243 227 245
rect 220 238 227 243
rect 233 240 238 247
rect 220 236 223 238
rect 225 236 227 238
rect 220 233 227 236
rect 231 238 238 240
rect 231 236 233 238
rect 235 236 238 238
rect 231 234 238 236
rect 200 230 205 233
rect 190 227 195 230
rect 233 227 238 234
rect 240 227 245 247
rect 247 241 254 247
rect 270 241 277 247
rect 279 245 287 247
rect 279 243 282 245
rect 284 243 287 245
rect 279 241 287 243
rect 289 241 297 247
rect 247 231 256 241
rect 247 229 250 231
rect 252 229 256 231
rect 247 227 256 229
rect 258 238 265 241
rect 258 236 261 238
rect 263 236 265 238
rect 258 234 265 236
rect 270 234 275 241
rect 291 238 297 241
rect 299 245 306 247
rect 299 243 302 245
rect 304 243 306 245
rect 299 241 306 243
rect 299 238 304 241
rect 384 244 392 246
rect 384 242 386 244
rect 388 242 392 244
rect 384 240 392 242
rect 394 244 402 246
rect 394 242 397 244
rect 399 242 402 244
rect 394 240 402 242
rect 404 244 411 246
rect 404 242 407 244
rect 409 242 411 244
rect 404 240 411 242
rect 607 241 614 243
rect 291 234 295 238
rect 258 227 263 234
rect 270 232 276 234
rect 270 230 272 232
rect 274 230 276 232
rect 270 228 276 230
rect 289 232 295 234
rect 314 237 321 239
rect 314 235 316 237
rect 318 235 321 237
rect 314 233 321 235
rect 323 237 331 239
rect 323 235 326 237
rect 328 235 331 237
rect 323 233 331 235
rect 333 233 338 239
rect 340 237 348 239
rect 340 235 343 237
rect 345 235 348 237
rect 340 233 348 235
rect 350 233 355 239
rect 357 237 365 239
rect 357 235 360 237
rect 362 235 365 237
rect 357 233 365 235
rect 367 237 374 239
rect 367 235 370 237
rect 372 235 374 237
rect 415 238 422 240
rect 415 236 417 238
rect 419 236 422 238
rect 367 233 374 235
rect 415 234 422 236
rect 424 238 432 240
rect 424 236 427 238
rect 429 236 432 238
rect 424 234 432 236
rect 434 234 439 240
rect 441 238 449 240
rect 441 236 444 238
rect 446 236 449 238
rect 441 234 449 236
rect 451 234 456 240
rect 458 238 466 240
rect 458 236 461 238
rect 463 236 466 238
rect 458 234 466 236
rect 468 238 475 240
rect 468 236 471 238
rect 473 236 475 238
rect 468 234 475 236
rect 479 238 486 240
rect 479 236 481 238
rect 483 236 486 238
rect 479 234 486 236
rect 488 238 496 240
rect 488 236 491 238
rect 493 236 496 238
rect 488 234 496 236
rect 498 234 503 240
rect 505 238 513 240
rect 505 236 508 238
rect 510 236 513 238
rect 505 234 513 236
rect 515 234 520 240
rect 522 238 530 240
rect 522 236 525 238
rect 527 236 530 238
rect 522 234 530 236
rect 532 238 539 240
rect 532 236 535 238
rect 537 236 539 238
rect 532 234 539 236
rect 543 238 550 240
rect 543 236 545 238
rect 547 236 550 238
rect 543 234 550 236
rect 552 238 560 240
rect 552 236 555 238
rect 557 236 560 238
rect 552 234 560 236
rect 562 234 567 240
rect 569 238 577 240
rect 569 236 572 238
rect 574 236 577 238
rect 569 234 577 236
rect 579 234 584 240
rect 586 238 594 240
rect 586 236 589 238
rect 591 236 594 238
rect 586 234 594 236
rect 596 238 603 240
rect 596 236 599 238
rect 601 236 603 238
rect 607 239 609 241
rect 611 239 614 241
rect 607 237 614 239
rect 616 241 624 243
rect 616 239 619 241
rect 621 239 624 241
rect 616 237 624 239
rect 626 241 634 243
rect 626 239 629 241
rect 631 239 634 241
rect 626 237 634 239
rect 636 241 643 243
rect 636 239 639 241
rect 641 239 643 241
rect 636 237 643 239
rect 648 241 655 243
rect 648 239 650 241
rect 652 239 655 241
rect 648 237 655 239
rect 657 240 665 243
rect 657 237 667 240
rect 596 234 603 236
rect 289 230 291 232
rect 293 230 295 232
rect 289 228 295 230
rect 659 231 667 237
rect 669 231 674 240
rect 676 238 683 240
rect 676 236 679 238
rect 681 236 683 238
rect 676 234 683 236
rect 676 231 681 234
rect 659 229 665 231
rect 659 227 661 229
rect 663 227 665 229
rect 659 225 665 227
rect 23 213 29 215
rect 23 211 25 213
rect 27 211 29 213
rect 23 209 29 211
rect 7 206 12 209
rect 5 204 12 206
rect 5 202 7 204
rect 9 202 12 204
rect 5 200 12 202
rect 14 200 19 209
rect 21 203 29 209
rect 393 210 399 212
rect 393 208 395 210
rect 397 208 399 210
rect 85 204 92 206
rect 21 200 31 203
rect 23 197 31 200
rect 33 201 40 203
rect 33 199 36 201
rect 38 199 40 201
rect 33 197 40 199
rect 45 201 52 203
rect 45 199 47 201
rect 49 199 52 201
rect 45 197 52 199
rect 54 201 62 203
rect 54 199 57 201
rect 59 199 62 201
rect 54 197 62 199
rect 64 201 72 203
rect 64 199 67 201
rect 69 199 72 201
rect 64 197 72 199
rect 74 201 81 203
rect 74 199 77 201
rect 79 199 81 201
rect 85 202 87 204
rect 89 202 92 204
rect 85 200 92 202
rect 94 204 102 206
rect 94 202 97 204
rect 99 202 102 204
rect 94 200 102 202
rect 104 200 109 206
rect 111 204 119 206
rect 111 202 114 204
rect 116 202 119 204
rect 111 200 119 202
rect 121 200 126 206
rect 128 204 136 206
rect 128 202 131 204
rect 133 202 136 204
rect 128 200 136 202
rect 138 204 145 206
rect 138 202 141 204
rect 143 202 145 204
rect 138 200 145 202
rect 149 204 156 206
rect 149 202 151 204
rect 153 202 156 204
rect 149 200 156 202
rect 158 204 166 206
rect 158 202 161 204
rect 163 202 166 204
rect 158 200 166 202
rect 168 200 173 206
rect 175 204 183 206
rect 175 202 178 204
rect 180 202 183 204
rect 175 200 183 202
rect 185 200 190 206
rect 192 204 200 206
rect 192 202 195 204
rect 197 202 200 204
rect 192 200 200 202
rect 202 204 209 206
rect 202 202 205 204
rect 207 202 209 204
rect 202 200 209 202
rect 213 204 220 206
rect 213 202 215 204
rect 217 202 220 204
rect 213 200 220 202
rect 222 204 230 206
rect 222 202 225 204
rect 227 202 230 204
rect 222 200 230 202
rect 232 200 237 206
rect 239 204 247 206
rect 239 202 242 204
rect 244 202 247 204
rect 239 200 247 202
rect 249 200 254 206
rect 256 204 264 206
rect 256 202 259 204
rect 261 202 264 204
rect 256 200 264 202
rect 266 204 273 206
rect 314 205 321 207
rect 266 202 269 204
rect 271 202 273 204
rect 266 200 273 202
rect 314 203 316 205
rect 318 203 321 205
rect 314 201 321 203
rect 323 205 331 207
rect 323 203 326 205
rect 328 203 331 205
rect 323 201 331 203
rect 333 201 338 207
rect 340 205 348 207
rect 340 203 343 205
rect 345 203 348 205
rect 340 201 348 203
rect 350 201 355 207
rect 357 205 365 207
rect 357 203 360 205
rect 362 203 365 205
rect 357 201 365 203
rect 367 205 374 207
rect 367 203 370 205
rect 372 203 374 205
rect 367 201 374 203
rect 393 206 399 208
rect 412 210 418 212
rect 412 208 414 210
rect 416 208 418 210
rect 412 206 418 208
rect 425 206 430 213
rect 393 202 397 206
rect 74 197 81 199
rect 277 198 284 200
rect 277 196 279 198
rect 281 196 284 198
rect 277 194 284 196
rect 286 198 294 200
rect 286 196 289 198
rect 291 196 294 198
rect 286 194 294 196
rect 296 198 304 200
rect 296 196 300 198
rect 302 196 304 198
rect 296 194 304 196
rect 384 199 389 202
rect 382 197 389 199
rect 382 195 384 197
rect 386 195 389 197
rect 382 193 389 195
rect 391 199 397 202
rect 413 199 418 206
rect 423 204 430 206
rect 423 202 425 204
rect 427 202 430 204
rect 423 199 430 202
rect 432 211 441 213
rect 432 209 436 211
rect 438 209 441 211
rect 432 199 441 209
rect 391 193 399 199
rect 401 197 409 199
rect 401 195 404 197
rect 406 195 409 197
rect 401 193 409 195
rect 411 193 418 199
rect 434 193 441 199
rect 443 193 448 213
rect 450 206 455 213
rect 493 210 498 213
rect 483 207 488 210
rect 450 204 457 206
rect 450 202 453 204
rect 455 202 457 204
rect 450 200 457 202
rect 461 204 468 207
rect 461 202 463 204
rect 465 202 468 204
rect 450 193 455 200
rect 461 197 468 202
rect 461 195 463 197
rect 465 195 468 197
rect 461 193 468 195
rect 470 197 478 207
rect 470 195 473 197
rect 475 195 478 197
rect 470 193 478 195
rect 480 205 488 207
rect 480 203 483 205
rect 485 203 488 205
rect 480 200 488 203
rect 490 208 498 210
rect 490 206 493 208
rect 495 206 498 208
rect 490 200 498 206
rect 500 206 505 213
rect 514 206 519 213
rect 500 204 507 206
rect 500 202 503 204
rect 505 202 507 204
rect 500 200 507 202
rect 512 204 519 206
rect 512 202 514 204
rect 516 202 519 204
rect 480 193 485 200
rect 512 199 519 202
rect 521 211 530 213
rect 521 209 525 211
rect 527 209 530 211
rect 521 199 530 209
rect 523 193 530 199
rect 532 193 537 213
rect 539 206 544 213
rect 582 210 587 213
rect 572 207 577 210
rect 539 204 546 206
rect 539 202 542 204
rect 544 202 546 204
rect 539 200 546 202
rect 550 204 557 207
rect 550 202 552 204
rect 554 202 557 204
rect 539 193 544 200
rect 550 197 557 202
rect 550 195 552 197
rect 554 195 557 197
rect 550 193 557 195
rect 559 197 567 207
rect 559 195 562 197
rect 564 195 567 197
rect 559 193 567 195
rect 569 205 577 207
rect 569 203 572 205
rect 574 203 577 205
rect 569 200 577 203
rect 579 208 587 210
rect 579 206 582 208
rect 584 206 587 208
rect 579 200 587 206
rect 589 206 594 213
rect 589 204 596 206
rect 611 205 617 207
rect 589 202 592 204
rect 594 202 596 204
rect 589 200 596 202
rect 600 203 607 205
rect 600 201 602 203
rect 604 201 607 203
rect 569 193 574 200
rect 600 199 607 201
rect 609 203 617 205
rect 609 201 612 203
rect 614 201 617 203
rect 609 199 617 201
rect 619 199 624 207
rect 626 205 634 207
rect 626 203 629 205
rect 631 203 634 205
rect 626 199 634 203
rect 636 199 641 207
rect 643 205 651 207
rect 643 203 646 205
rect 648 203 651 205
rect 643 199 651 203
rect 646 198 651 199
rect 653 204 658 207
rect 653 202 660 204
rect 653 200 656 202
rect 658 200 660 202
rect 653 198 660 200
rect 666 199 671 202
rect 664 197 671 199
rect 664 195 666 197
rect 668 195 671 197
rect 664 193 671 195
rect 673 200 684 202
rect 673 198 680 200
rect 682 198 684 200
rect 673 193 684 198
rect 4 95 15 100
rect 4 93 6 95
rect 8 93 15 95
rect 4 91 15 93
rect 17 98 24 100
rect 17 96 20 98
rect 22 96 24 98
rect 17 94 24 96
rect 17 91 22 94
rect 28 93 35 95
rect 28 91 30 93
rect 32 91 35 93
rect 28 89 35 91
rect 30 86 35 89
rect 37 94 42 95
rect 37 90 45 94
rect 37 88 40 90
rect 42 88 45 90
rect 37 86 45 88
rect 47 86 52 94
rect 54 90 62 94
rect 54 88 57 90
rect 59 88 62 90
rect 54 86 62 88
rect 64 86 69 94
rect 71 92 79 94
rect 71 90 74 92
rect 76 90 79 92
rect 71 88 79 90
rect 81 92 88 94
rect 114 93 119 100
rect 81 90 84 92
rect 86 90 88 92
rect 81 88 88 90
rect 92 91 99 93
rect 92 89 94 91
rect 96 89 99 91
rect 71 86 77 88
rect 92 87 99 89
rect 94 80 99 87
rect 101 87 109 93
rect 101 85 104 87
rect 106 85 109 87
rect 101 83 109 85
rect 111 90 119 93
rect 111 88 114 90
rect 116 88 119 90
rect 111 86 119 88
rect 121 98 129 100
rect 121 96 124 98
rect 126 96 129 98
rect 121 86 129 96
rect 131 98 138 100
rect 131 96 134 98
rect 136 96 138 98
rect 131 91 138 96
rect 144 93 149 100
rect 131 89 134 91
rect 136 89 138 91
rect 131 86 138 89
rect 142 91 149 93
rect 142 89 144 91
rect 146 89 149 91
rect 142 87 149 89
rect 111 83 116 86
rect 101 80 106 83
rect 144 80 149 87
rect 151 80 156 100
rect 158 94 165 100
rect 158 84 167 94
rect 158 82 161 84
rect 163 82 167 84
rect 158 80 167 82
rect 169 91 176 94
rect 203 93 208 100
rect 169 89 172 91
rect 174 89 176 91
rect 169 87 176 89
rect 181 91 188 93
rect 181 89 183 91
rect 185 89 188 91
rect 181 87 188 89
rect 169 80 174 87
rect 183 80 188 87
rect 190 87 198 93
rect 190 85 193 87
rect 195 85 198 87
rect 190 83 198 85
rect 200 90 208 93
rect 200 88 203 90
rect 205 88 208 90
rect 200 86 208 88
rect 210 98 218 100
rect 210 96 213 98
rect 215 96 218 98
rect 210 86 218 96
rect 220 98 227 100
rect 220 96 223 98
rect 225 96 227 98
rect 220 91 227 96
rect 233 93 238 100
rect 220 89 223 91
rect 225 89 227 91
rect 220 86 227 89
rect 231 91 238 93
rect 231 89 233 91
rect 235 89 238 91
rect 231 87 238 89
rect 200 83 205 86
rect 190 80 195 83
rect 233 80 238 87
rect 240 80 245 100
rect 247 94 254 100
rect 270 94 277 100
rect 279 98 287 100
rect 279 96 282 98
rect 284 96 287 98
rect 279 94 287 96
rect 289 94 297 100
rect 247 84 256 94
rect 247 82 250 84
rect 252 82 256 84
rect 247 80 256 82
rect 258 91 265 94
rect 258 89 261 91
rect 263 89 265 91
rect 258 87 265 89
rect 270 87 275 94
rect 291 91 297 94
rect 299 98 306 100
rect 299 96 302 98
rect 304 96 306 98
rect 299 94 306 96
rect 299 91 304 94
rect 384 97 392 99
rect 384 95 386 97
rect 388 95 392 97
rect 384 93 392 95
rect 394 97 402 99
rect 394 95 397 97
rect 399 95 402 97
rect 394 93 402 95
rect 404 97 411 99
rect 404 95 407 97
rect 409 95 411 97
rect 404 93 411 95
rect 607 94 614 96
rect 291 87 295 91
rect 258 80 263 87
rect 270 85 276 87
rect 270 83 272 85
rect 274 83 276 85
rect 270 81 276 83
rect 289 85 295 87
rect 314 90 321 92
rect 314 88 316 90
rect 318 88 321 90
rect 314 86 321 88
rect 323 90 331 92
rect 323 88 326 90
rect 328 88 331 90
rect 323 86 331 88
rect 333 86 338 92
rect 340 90 348 92
rect 340 88 343 90
rect 345 88 348 90
rect 340 86 348 88
rect 350 86 355 92
rect 357 90 365 92
rect 357 88 360 90
rect 362 88 365 90
rect 357 86 365 88
rect 367 90 374 92
rect 367 88 370 90
rect 372 88 374 90
rect 415 91 422 93
rect 415 89 417 91
rect 419 89 422 91
rect 367 86 374 88
rect 415 87 422 89
rect 424 91 432 93
rect 424 89 427 91
rect 429 89 432 91
rect 424 87 432 89
rect 434 87 439 93
rect 441 91 449 93
rect 441 89 444 91
rect 446 89 449 91
rect 441 87 449 89
rect 451 87 456 93
rect 458 91 466 93
rect 458 89 461 91
rect 463 89 466 91
rect 458 87 466 89
rect 468 91 475 93
rect 468 89 471 91
rect 473 89 475 91
rect 468 87 475 89
rect 479 91 486 93
rect 479 89 481 91
rect 483 89 486 91
rect 479 87 486 89
rect 488 91 496 93
rect 488 89 491 91
rect 493 89 496 91
rect 488 87 496 89
rect 498 87 503 93
rect 505 91 513 93
rect 505 89 508 91
rect 510 89 513 91
rect 505 87 513 89
rect 515 87 520 93
rect 522 91 530 93
rect 522 89 525 91
rect 527 89 530 91
rect 522 87 530 89
rect 532 91 539 93
rect 532 89 535 91
rect 537 89 539 91
rect 532 87 539 89
rect 543 91 550 93
rect 543 89 545 91
rect 547 89 550 91
rect 543 87 550 89
rect 552 91 560 93
rect 552 89 555 91
rect 557 89 560 91
rect 552 87 560 89
rect 562 87 567 93
rect 569 91 577 93
rect 569 89 572 91
rect 574 89 577 91
rect 569 87 577 89
rect 579 87 584 93
rect 586 91 594 93
rect 586 89 589 91
rect 591 89 594 91
rect 586 87 594 89
rect 596 91 603 93
rect 596 89 599 91
rect 601 89 603 91
rect 607 92 609 94
rect 611 92 614 94
rect 607 90 614 92
rect 616 94 624 96
rect 616 92 619 94
rect 621 92 624 94
rect 616 90 624 92
rect 626 94 634 96
rect 626 92 629 94
rect 631 92 634 94
rect 626 90 634 92
rect 636 94 643 96
rect 636 92 639 94
rect 641 92 643 94
rect 636 90 643 92
rect 648 94 655 96
rect 648 92 650 94
rect 652 92 655 94
rect 648 90 655 92
rect 657 93 665 96
rect 657 90 667 93
rect 596 87 603 89
rect 289 83 291 85
rect 293 83 295 85
rect 289 81 295 83
rect 659 84 667 90
rect 669 84 674 93
rect 676 91 683 93
rect 676 89 679 91
rect 681 89 683 91
rect 676 87 683 89
rect 676 84 681 87
rect 659 82 665 84
rect 659 80 661 82
rect 663 80 665 82
rect 659 78 665 80
rect 23 66 29 68
rect 23 64 25 66
rect 27 64 29 66
rect 23 62 29 64
rect 7 59 12 62
rect 5 57 12 59
rect 5 55 7 57
rect 9 55 12 57
rect 5 53 12 55
rect 14 53 19 62
rect 21 56 29 62
rect 393 63 399 65
rect 393 61 395 63
rect 397 61 399 63
rect 85 57 92 59
rect 21 53 31 56
rect 23 50 31 53
rect 33 54 40 56
rect 33 52 36 54
rect 38 52 40 54
rect 33 50 40 52
rect 45 54 52 56
rect 45 52 47 54
rect 49 52 52 54
rect 45 50 52 52
rect 54 54 62 56
rect 54 52 57 54
rect 59 52 62 54
rect 54 50 62 52
rect 64 54 72 56
rect 64 52 67 54
rect 69 52 72 54
rect 64 50 72 52
rect 74 54 81 56
rect 74 52 77 54
rect 79 52 81 54
rect 85 55 87 57
rect 89 55 92 57
rect 85 53 92 55
rect 94 57 102 59
rect 94 55 97 57
rect 99 55 102 57
rect 94 53 102 55
rect 104 53 109 59
rect 111 57 119 59
rect 111 55 114 57
rect 116 55 119 57
rect 111 53 119 55
rect 121 53 126 59
rect 128 57 136 59
rect 128 55 131 57
rect 133 55 136 57
rect 128 53 136 55
rect 138 57 145 59
rect 138 55 141 57
rect 143 55 145 57
rect 138 53 145 55
rect 149 57 156 59
rect 149 55 151 57
rect 153 55 156 57
rect 149 53 156 55
rect 158 57 166 59
rect 158 55 161 57
rect 163 55 166 57
rect 158 53 166 55
rect 168 53 173 59
rect 175 57 183 59
rect 175 55 178 57
rect 180 55 183 57
rect 175 53 183 55
rect 185 53 190 59
rect 192 57 200 59
rect 192 55 195 57
rect 197 55 200 57
rect 192 53 200 55
rect 202 57 209 59
rect 202 55 205 57
rect 207 55 209 57
rect 202 53 209 55
rect 213 57 220 59
rect 213 55 215 57
rect 217 55 220 57
rect 213 53 220 55
rect 222 57 230 59
rect 222 55 225 57
rect 227 55 230 57
rect 222 53 230 55
rect 232 53 237 59
rect 239 57 247 59
rect 239 55 242 57
rect 244 55 247 57
rect 239 53 247 55
rect 249 53 254 59
rect 256 57 264 59
rect 256 55 259 57
rect 261 55 264 57
rect 256 53 264 55
rect 266 57 273 59
rect 314 58 321 60
rect 266 55 269 57
rect 271 55 273 57
rect 266 53 273 55
rect 314 56 316 58
rect 318 56 321 58
rect 314 54 321 56
rect 323 58 331 60
rect 323 56 326 58
rect 328 56 331 58
rect 323 54 331 56
rect 333 54 338 60
rect 340 58 348 60
rect 340 56 343 58
rect 345 56 348 58
rect 340 54 348 56
rect 350 54 355 60
rect 357 58 365 60
rect 357 56 360 58
rect 362 56 365 58
rect 357 54 365 56
rect 367 58 374 60
rect 367 56 370 58
rect 372 56 374 58
rect 367 54 374 56
rect 393 59 399 61
rect 412 63 418 65
rect 412 61 414 63
rect 416 61 418 63
rect 412 59 418 61
rect 425 59 430 66
rect 393 55 397 59
rect 74 50 81 52
rect 277 51 284 53
rect 277 49 279 51
rect 281 49 284 51
rect 277 47 284 49
rect 286 51 294 53
rect 286 49 289 51
rect 291 49 294 51
rect 286 47 294 49
rect 296 51 304 53
rect 296 49 300 51
rect 302 49 304 51
rect 296 47 304 49
rect 384 52 389 55
rect 382 50 389 52
rect 382 48 384 50
rect 386 48 389 50
rect 382 46 389 48
rect 391 52 397 55
rect 413 52 418 59
rect 423 57 430 59
rect 423 55 425 57
rect 427 55 430 57
rect 423 52 430 55
rect 432 64 441 66
rect 432 62 436 64
rect 438 62 441 64
rect 432 52 441 62
rect 391 46 399 52
rect 401 50 409 52
rect 401 48 404 50
rect 406 48 409 50
rect 401 46 409 48
rect 411 46 418 52
rect 434 46 441 52
rect 443 46 448 66
rect 450 59 455 66
rect 493 63 498 66
rect 483 60 488 63
rect 450 57 457 59
rect 450 55 453 57
rect 455 55 457 57
rect 450 53 457 55
rect 461 57 468 60
rect 461 55 463 57
rect 465 55 468 57
rect 450 46 455 53
rect 461 50 468 55
rect 461 48 463 50
rect 465 48 468 50
rect 461 46 468 48
rect 470 50 478 60
rect 470 48 473 50
rect 475 48 478 50
rect 470 46 478 48
rect 480 58 488 60
rect 480 56 483 58
rect 485 56 488 58
rect 480 53 488 56
rect 490 61 498 63
rect 490 59 493 61
rect 495 59 498 61
rect 490 53 498 59
rect 500 59 505 66
rect 514 59 519 66
rect 500 57 507 59
rect 500 55 503 57
rect 505 55 507 57
rect 500 53 507 55
rect 512 57 519 59
rect 512 55 514 57
rect 516 55 519 57
rect 480 46 485 53
rect 512 52 519 55
rect 521 64 530 66
rect 521 62 525 64
rect 527 62 530 64
rect 521 52 530 62
rect 523 46 530 52
rect 532 46 537 66
rect 539 59 544 66
rect 582 63 587 66
rect 572 60 577 63
rect 539 57 546 59
rect 539 55 542 57
rect 544 55 546 57
rect 539 53 546 55
rect 550 57 557 60
rect 550 55 552 57
rect 554 55 557 57
rect 539 46 544 53
rect 550 50 557 55
rect 550 48 552 50
rect 554 48 557 50
rect 550 46 557 48
rect 559 50 567 60
rect 559 48 562 50
rect 564 48 567 50
rect 559 46 567 48
rect 569 58 577 60
rect 569 56 572 58
rect 574 56 577 58
rect 569 53 577 56
rect 579 61 587 63
rect 579 59 582 61
rect 584 59 587 61
rect 579 53 587 59
rect 589 59 594 66
rect 589 57 596 59
rect 611 58 617 60
rect 589 55 592 57
rect 594 55 596 57
rect 589 53 596 55
rect 600 56 607 58
rect 600 54 602 56
rect 604 54 607 56
rect 569 46 574 53
rect 600 52 607 54
rect 609 56 617 58
rect 609 54 612 56
rect 614 54 617 56
rect 609 52 617 54
rect 619 52 624 60
rect 626 58 634 60
rect 626 56 629 58
rect 631 56 634 58
rect 626 52 634 56
rect 636 52 641 60
rect 643 58 651 60
rect 643 56 646 58
rect 648 56 651 58
rect 643 52 651 56
rect 646 51 651 52
rect 653 57 658 60
rect 653 55 660 57
rect 653 53 656 55
rect 658 53 660 55
rect 653 51 660 53
rect 666 52 671 55
rect 664 50 671 52
rect 664 48 666 50
rect 668 48 671 50
rect 664 46 671 48
rect 673 53 684 55
rect 673 51 680 53
rect 682 51 684 53
rect 673 46 684 51
<< pdif >>
rect 6 278 13 280
rect 6 276 9 278
rect 11 277 13 278
rect 30 280 35 287
rect 28 278 35 280
rect 11 276 15 277
rect 6 259 15 276
rect 17 272 22 277
rect 28 276 30 278
rect 32 276 35 278
rect 28 274 35 276
rect 17 270 24 272
rect 17 268 20 270
rect 22 268 24 270
rect 30 269 35 274
rect 37 285 45 287
rect 37 283 40 285
rect 42 283 45 285
rect 37 271 45 283
rect 47 271 52 287
rect 54 275 62 287
rect 54 273 57 275
rect 59 273 62 275
rect 54 271 62 273
rect 64 271 69 287
rect 71 285 78 287
rect 71 283 74 285
rect 76 283 78 285
rect 71 275 78 283
rect 71 271 77 275
rect 94 275 99 287
rect 37 269 42 271
rect 17 263 24 268
rect 17 261 20 263
rect 22 261 24 263
rect 17 259 24 261
rect 73 267 77 271
rect 92 273 99 275
rect 92 271 94 273
rect 96 271 99 273
rect 73 259 79 267
rect 81 265 86 267
rect 92 266 99 271
rect 81 263 88 265
rect 81 261 84 263
rect 86 261 88 263
rect 92 264 94 266
rect 96 264 99 266
rect 92 262 99 264
rect 101 285 110 287
rect 101 283 105 285
rect 107 283 110 285
rect 133 285 147 287
rect 133 284 140 285
rect 101 275 110 283
rect 117 275 122 284
rect 101 262 112 275
rect 114 266 122 275
rect 114 264 117 266
rect 119 264 122 266
rect 114 262 122 264
rect 81 259 88 261
rect 117 259 122 262
rect 124 259 129 284
rect 131 283 140 284
rect 142 283 147 285
rect 131 278 147 283
rect 131 276 140 278
rect 142 276 147 278
rect 131 259 147 276
rect 149 277 157 287
rect 149 275 152 277
rect 154 275 157 277
rect 149 270 157 275
rect 149 268 152 270
rect 154 268 157 270
rect 149 259 157 268
rect 159 285 167 287
rect 159 283 162 285
rect 164 283 167 285
rect 159 278 167 283
rect 159 276 162 278
rect 164 276 167 278
rect 159 259 167 276
rect 169 272 174 287
rect 183 275 188 287
rect 181 273 188 275
rect 169 270 176 272
rect 169 268 172 270
rect 174 268 176 270
rect 169 263 176 268
rect 169 261 172 263
rect 174 261 176 263
rect 181 271 183 273
rect 185 271 188 273
rect 181 266 188 271
rect 181 264 183 266
rect 185 264 188 266
rect 181 262 188 264
rect 190 285 199 287
rect 190 283 194 285
rect 196 283 199 285
rect 222 285 236 287
rect 222 284 229 285
rect 190 275 199 283
rect 206 275 211 284
rect 190 262 201 275
rect 203 266 211 275
rect 203 264 206 266
rect 208 264 211 266
rect 203 262 211 264
rect 169 259 176 261
rect 206 259 211 262
rect 213 259 218 284
rect 220 283 229 284
rect 231 283 236 285
rect 220 278 236 283
rect 220 276 229 278
rect 231 276 236 278
rect 220 259 236 276
rect 238 277 246 287
rect 238 275 241 277
rect 243 275 246 277
rect 238 270 246 275
rect 238 268 241 270
rect 243 268 246 270
rect 238 259 246 268
rect 248 285 256 287
rect 248 283 251 285
rect 253 283 256 285
rect 248 278 256 283
rect 248 276 251 278
rect 253 276 256 278
rect 248 259 256 276
rect 258 272 263 287
rect 272 280 277 287
rect 270 278 277 280
rect 270 276 272 278
rect 274 276 277 278
rect 270 274 277 276
rect 258 270 265 272
rect 258 268 261 270
rect 263 268 265 270
rect 258 263 265 268
rect 272 266 277 274
rect 279 266 284 287
rect 286 285 295 287
rect 286 283 291 285
rect 293 283 295 285
rect 286 277 295 283
rect 389 281 394 287
rect 387 279 394 281
rect 286 266 297 277
rect 258 261 261 263
rect 263 261 265 263
rect 258 259 265 261
rect 289 259 297 266
rect 299 275 306 277
rect 299 273 302 275
rect 304 273 306 275
rect 316 273 321 279
rect 299 268 306 273
rect 299 266 302 268
rect 304 266 306 268
rect 314 271 321 273
rect 314 269 316 271
rect 318 269 321 271
rect 314 267 321 269
rect 323 277 331 279
rect 323 275 326 277
rect 328 275 331 277
rect 323 267 331 275
rect 333 267 338 279
rect 340 271 348 279
rect 340 269 343 271
rect 345 269 348 271
rect 340 267 348 269
rect 350 267 355 279
rect 357 277 364 279
rect 357 275 360 277
rect 362 275 364 277
rect 387 277 389 279
rect 391 277 394 279
rect 387 275 394 277
rect 357 273 364 275
rect 357 267 363 273
rect 299 264 306 266
rect 299 259 304 264
rect 359 265 363 267
rect 389 267 394 275
rect 396 267 401 287
rect 403 285 412 287
rect 618 286 627 288
rect 403 283 408 285
rect 410 283 412 285
rect 403 278 412 283
rect 618 284 621 286
rect 623 284 627 286
rect 403 276 408 278
rect 410 276 412 278
rect 403 273 412 276
rect 425 278 432 280
rect 425 276 427 278
rect 429 276 432 278
rect 425 274 432 276
rect 403 267 411 273
rect 359 259 365 265
rect 367 263 374 265
rect 367 261 370 263
rect 372 261 374 263
rect 367 259 374 261
rect 426 268 432 274
rect 434 268 439 280
rect 441 272 449 280
rect 441 270 444 272
rect 446 270 449 272
rect 441 268 449 270
rect 451 268 456 280
rect 458 278 466 280
rect 458 276 461 278
rect 463 276 466 278
rect 458 268 466 276
rect 468 274 473 280
rect 481 274 486 280
rect 468 272 475 274
rect 468 270 471 272
rect 473 270 475 272
rect 468 268 475 270
rect 479 272 486 274
rect 479 270 481 272
rect 483 270 486 272
rect 479 268 486 270
rect 488 278 496 280
rect 488 276 491 278
rect 493 276 496 278
rect 488 268 496 276
rect 498 268 503 280
rect 505 272 513 280
rect 505 270 508 272
rect 510 270 513 272
rect 505 268 513 270
rect 515 268 520 280
rect 522 278 529 280
rect 522 276 525 278
rect 527 276 529 278
rect 522 274 529 276
rect 522 268 528 274
rect 545 274 550 280
rect 426 266 430 268
rect 415 264 422 266
rect 415 262 417 264
rect 419 262 422 264
rect 415 260 422 262
rect 424 260 430 266
rect 524 266 528 268
rect 543 272 550 274
rect 543 270 545 272
rect 547 270 550 272
rect 543 268 550 270
rect 552 278 560 280
rect 552 276 555 278
rect 557 276 560 278
rect 552 268 560 276
rect 562 268 567 280
rect 569 272 577 280
rect 569 270 572 272
rect 574 270 577 272
rect 569 268 577 270
rect 579 268 584 280
rect 586 278 593 280
rect 618 279 627 284
rect 586 276 589 278
rect 591 276 593 278
rect 586 274 593 276
rect 607 277 614 279
rect 607 275 609 277
rect 611 275 614 277
rect 586 268 592 274
rect 607 273 614 275
rect 524 260 530 266
rect 532 264 539 266
rect 532 262 535 264
rect 537 262 539 264
rect 532 260 539 262
rect 588 266 592 268
rect 609 267 614 273
rect 616 270 627 279
rect 629 270 634 288
rect 636 281 641 288
rect 636 279 643 281
rect 636 277 639 279
rect 641 277 643 279
rect 636 275 643 277
rect 636 270 641 275
rect 616 267 624 270
rect 588 260 594 266
rect 596 264 603 266
rect 596 262 599 264
rect 601 262 603 264
rect 596 260 603 262
rect 650 266 655 272
rect 648 264 655 266
rect 648 262 650 264
rect 652 262 655 264
rect 648 260 655 262
rect 657 270 663 272
rect 657 264 665 270
rect 657 262 660 264
rect 662 262 665 264
rect 657 260 665 262
rect 667 264 675 270
rect 667 262 670 264
rect 672 262 675 264
rect 667 260 675 262
rect 677 268 684 270
rect 677 266 680 268
rect 682 266 684 268
rect 677 260 684 266
rect 4 174 11 180
rect 4 172 6 174
rect 8 172 11 174
rect 4 170 11 172
rect 13 178 21 180
rect 13 176 16 178
rect 18 176 21 178
rect 13 170 21 176
rect 23 178 31 180
rect 23 176 26 178
rect 28 176 31 178
rect 23 170 31 176
rect 25 168 31 170
rect 33 178 40 180
rect 33 176 36 178
rect 38 176 40 178
rect 33 174 40 176
rect 33 168 38 174
rect 85 178 92 180
rect 85 176 87 178
rect 89 176 92 178
rect 85 174 92 176
rect 94 174 100 180
rect 64 170 72 173
rect 47 165 52 170
rect 45 163 52 165
rect 45 161 47 163
rect 49 161 52 163
rect 45 159 52 161
rect 47 152 52 159
rect 54 152 59 170
rect 61 161 72 170
rect 74 167 79 173
rect 96 172 100 174
rect 149 178 156 180
rect 149 176 151 178
rect 153 176 156 178
rect 149 174 156 176
rect 158 174 164 180
rect 74 165 81 167
rect 96 166 102 172
rect 74 163 77 165
rect 79 163 81 165
rect 74 161 81 163
rect 95 164 102 166
rect 95 162 97 164
rect 99 162 102 164
rect 61 156 70 161
rect 95 160 102 162
rect 104 160 109 172
rect 111 170 119 172
rect 111 168 114 170
rect 116 168 119 170
rect 111 160 119 168
rect 121 160 126 172
rect 128 164 136 172
rect 128 162 131 164
rect 133 162 136 164
rect 128 160 136 162
rect 138 170 145 172
rect 138 168 141 170
rect 143 168 145 170
rect 138 166 145 168
rect 160 172 164 174
rect 258 174 264 180
rect 266 178 273 180
rect 266 176 269 178
rect 271 176 273 178
rect 266 174 273 176
rect 258 172 262 174
rect 138 160 143 166
rect 160 166 166 172
rect 159 164 166 166
rect 159 162 161 164
rect 163 162 166 164
rect 159 160 166 162
rect 168 160 173 172
rect 175 170 183 172
rect 175 168 178 170
rect 180 168 183 170
rect 175 160 183 168
rect 185 160 190 172
rect 192 164 200 172
rect 192 162 195 164
rect 197 162 200 164
rect 192 160 200 162
rect 202 170 209 172
rect 202 168 205 170
rect 207 168 209 170
rect 202 166 209 168
rect 213 170 220 172
rect 213 168 215 170
rect 217 168 220 170
rect 213 166 220 168
rect 202 160 207 166
rect 215 160 220 166
rect 222 164 230 172
rect 222 162 225 164
rect 227 162 230 164
rect 222 160 230 162
rect 232 160 237 172
rect 239 170 247 172
rect 239 168 242 170
rect 244 168 247 170
rect 239 160 247 168
rect 249 160 254 172
rect 256 166 262 172
rect 314 179 321 181
rect 314 177 316 179
rect 318 177 321 179
rect 314 175 321 177
rect 323 175 329 181
rect 277 167 285 173
rect 256 164 263 166
rect 256 162 259 164
rect 261 162 263 164
rect 256 160 263 162
rect 276 164 285 167
rect 276 162 278 164
rect 280 162 285 164
rect 61 154 65 156
rect 67 154 70 156
rect 276 157 285 162
rect 276 155 278 157
rect 280 155 285 157
rect 61 152 70 154
rect 276 153 285 155
rect 287 153 292 173
rect 294 165 299 173
rect 325 173 329 175
rect 384 176 389 181
rect 382 174 389 176
rect 325 167 331 173
rect 324 165 331 167
rect 294 163 301 165
rect 294 161 297 163
rect 299 161 301 163
rect 324 163 326 165
rect 328 163 331 165
rect 324 161 331 163
rect 333 161 338 173
rect 340 171 348 173
rect 340 169 343 171
rect 345 169 348 171
rect 340 161 348 169
rect 350 161 355 173
rect 357 165 365 173
rect 357 163 360 165
rect 362 163 365 165
rect 357 161 365 163
rect 367 171 374 173
rect 367 169 370 171
rect 372 169 374 171
rect 367 167 374 169
rect 382 172 384 174
rect 386 172 389 174
rect 382 167 389 172
rect 367 161 372 167
rect 382 165 384 167
rect 386 165 389 167
rect 382 163 389 165
rect 391 174 399 181
rect 423 179 430 181
rect 423 177 425 179
rect 427 177 430 179
rect 391 163 402 174
rect 294 159 301 161
rect 294 153 299 159
rect 393 157 402 163
rect 393 155 395 157
rect 397 155 402 157
rect 393 153 402 155
rect 404 153 409 174
rect 411 166 416 174
rect 423 172 430 177
rect 423 170 425 172
rect 427 170 430 172
rect 423 168 430 170
rect 411 164 418 166
rect 411 162 414 164
rect 416 162 418 164
rect 411 160 418 162
rect 411 153 416 160
rect 425 153 430 168
rect 432 164 440 181
rect 432 162 435 164
rect 437 162 440 164
rect 432 157 440 162
rect 432 155 435 157
rect 437 155 440 157
rect 432 153 440 155
rect 442 172 450 181
rect 442 170 445 172
rect 447 170 450 172
rect 442 165 450 170
rect 442 163 445 165
rect 447 163 450 165
rect 442 153 450 163
rect 452 164 468 181
rect 452 162 457 164
rect 459 162 468 164
rect 452 157 468 162
rect 452 155 457 157
rect 459 156 468 157
rect 470 156 475 181
rect 477 178 482 181
rect 512 179 519 181
rect 477 176 485 178
rect 477 174 480 176
rect 482 174 485 176
rect 477 165 485 174
rect 487 165 498 178
rect 477 156 482 165
rect 489 157 498 165
rect 459 155 466 156
rect 452 153 466 155
rect 489 155 492 157
rect 494 155 498 157
rect 489 153 498 155
rect 500 176 507 178
rect 500 174 503 176
rect 505 174 507 176
rect 500 169 507 174
rect 500 167 503 169
rect 505 167 507 169
rect 512 177 514 179
rect 516 177 519 179
rect 512 172 519 177
rect 512 170 514 172
rect 516 170 519 172
rect 512 168 519 170
rect 500 165 507 167
rect 500 153 505 165
rect 514 153 519 168
rect 521 164 529 181
rect 521 162 524 164
rect 526 162 529 164
rect 521 157 529 162
rect 521 155 524 157
rect 526 155 529 157
rect 521 153 529 155
rect 531 172 539 181
rect 531 170 534 172
rect 536 170 539 172
rect 531 165 539 170
rect 531 163 534 165
rect 536 163 539 165
rect 531 153 539 163
rect 541 164 557 181
rect 541 162 546 164
rect 548 162 557 164
rect 541 157 557 162
rect 541 155 546 157
rect 548 156 557 157
rect 559 156 564 181
rect 566 178 571 181
rect 600 179 607 181
rect 566 176 574 178
rect 566 174 569 176
rect 571 174 574 176
rect 566 165 574 174
rect 576 165 587 178
rect 566 156 571 165
rect 578 157 587 165
rect 548 155 555 156
rect 541 153 555 155
rect 578 155 581 157
rect 583 155 587 157
rect 578 153 587 155
rect 589 176 596 178
rect 589 174 592 176
rect 594 174 596 176
rect 600 177 602 179
rect 604 177 607 179
rect 600 175 607 177
rect 589 169 596 174
rect 602 173 607 175
rect 609 173 615 181
rect 589 167 592 169
rect 594 167 596 169
rect 589 165 596 167
rect 611 169 615 173
rect 664 179 671 181
rect 664 177 666 179
rect 668 177 671 179
rect 664 172 671 177
rect 646 169 651 171
rect 589 153 594 165
rect 611 165 617 169
rect 610 157 617 165
rect 610 155 612 157
rect 614 155 617 157
rect 610 153 617 155
rect 619 153 624 169
rect 626 167 634 169
rect 626 165 629 167
rect 631 165 634 167
rect 626 153 634 165
rect 636 153 641 169
rect 643 157 651 169
rect 643 155 646 157
rect 648 155 651 157
rect 643 153 651 155
rect 653 166 658 171
rect 664 170 666 172
rect 668 170 671 172
rect 664 168 671 170
rect 653 164 660 166
rect 653 162 656 164
rect 658 162 660 164
rect 666 163 671 168
rect 673 164 682 181
rect 673 163 677 164
rect 653 160 660 162
rect 653 153 658 160
rect 675 162 677 163
rect 679 162 682 164
rect 675 160 682 162
rect 6 131 13 133
rect 6 129 9 131
rect 11 130 13 131
rect 30 133 35 140
rect 28 131 35 133
rect 11 129 15 130
rect 6 112 15 129
rect 17 125 22 130
rect 28 129 30 131
rect 32 129 35 131
rect 28 127 35 129
rect 17 123 24 125
rect 17 121 20 123
rect 22 121 24 123
rect 30 122 35 127
rect 37 138 45 140
rect 37 136 40 138
rect 42 136 45 138
rect 37 124 45 136
rect 47 124 52 140
rect 54 128 62 140
rect 54 126 57 128
rect 59 126 62 128
rect 54 124 62 126
rect 64 124 69 140
rect 71 138 78 140
rect 71 136 74 138
rect 76 136 78 138
rect 71 128 78 136
rect 71 124 77 128
rect 94 128 99 140
rect 37 122 42 124
rect 17 116 24 121
rect 17 114 20 116
rect 22 114 24 116
rect 17 112 24 114
rect 73 120 77 124
rect 92 126 99 128
rect 92 124 94 126
rect 96 124 99 126
rect 73 112 79 120
rect 81 118 86 120
rect 92 119 99 124
rect 81 116 88 118
rect 81 114 84 116
rect 86 114 88 116
rect 92 117 94 119
rect 96 117 99 119
rect 92 115 99 117
rect 101 138 110 140
rect 101 136 105 138
rect 107 136 110 138
rect 133 138 147 140
rect 133 137 140 138
rect 101 128 110 136
rect 117 128 122 137
rect 101 115 112 128
rect 114 119 122 128
rect 114 117 117 119
rect 119 117 122 119
rect 114 115 122 117
rect 81 112 88 114
rect 117 112 122 115
rect 124 112 129 137
rect 131 136 140 137
rect 142 136 147 138
rect 131 131 147 136
rect 131 129 140 131
rect 142 129 147 131
rect 131 112 147 129
rect 149 130 157 140
rect 149 128 152 130
rect 154 128 157 130
rect 149 123 157 128
rect 149 121 152 123
rect 154 121 157 123
rect 149 112 157 121
rect 159 138 167 140
rect 159 136 162 138
rect 164 136 167 138
rect 159 131 167 136
rect 159 129 162 131
rect 164 129 167 131
rect 159 112 167 129
rect 169 125 174 140
rect 183 128 188 140
rect 181 126 188 128
rect 169 123 176 125
rect 169 121 172 123
rect 174 121 176 123
rect 169 116 176 121
rect 169 114 172 116
rect 174 114 176 116
rect 181 124 183 126
rect 185 124 188 126
rect 181 119 188 124
rect 181 117 183 119
rect 185 117 188 119
rect 181 115 188 117
rect 190 138 199 140
rect 190 136 194 138
rect 196 136 199 138
rect 222 138 236 140
rect 222 137 229 138
rect 190 128 199 136
rect 206 128 211 137
rect 190 115 201 128
rect 203 119 211 128
rect 203 117 206 119
rect 208 117 211 119
rect 203 115 211 117
rect 169 112 176 114
rect 206 112 211 115
rect 213 112 218 137
rect 220 136 229 137
rect 231 136 236 138
rect 220 131 236 136
rect 220 129 229 131
rect 231 129 236 131
rect 220 112 236 129
rect 238 130 246 140
rect 238 128 241 130
rect 243 128 246 130
rect 238 123 246 128
rect 238 121 241 123
rect 243 121 246 123
rect 238 112 246 121
rect 248 138 256 140
rect 248 136 251 138
rect 253 136 256 138
rect 248 131 256 136
rect 248 129 251 131
rect 253 129 256 131
rect 248 112 256 129
rect 258 125 263 140
rect 272 133 277 140
rect 270 131 277 133
rect 270 129 272 131
rect 274 129 277 131
rect 270 127 277 129
rect 258 123 265 125
rect 258 121 261 123
rect 263 121 265 123
rect 258 116 265 121
rect 272 119 277 127
rect 279 119 284 140
rect 286 138 295 140
rect 286 136 291 138
rect 293 136 295 138
rect 286 130 295 136
rect 389 134 394 140
rect 387 132 394 134
rect 286 119 297 130
rect 258 114 261 116
rect 263 114 265 116
rect 258 112 265 114
rect 289 112 297 119
rect 299 128 306 130
rect 299 126 302 128
rect 304 126 306 128
rect 316 126 321 132
rect 299 121 306 126
rect 299 119 302 121
rect 304 119 306 121
rect 314 124 321 126
rect 314 122 316 124
rect 318 122 321 124
rect 314 120 321 122
rect 323 130 331 132
rect 323 128 326 130
rect 328 128 331 130
rect 323 120 331 128
rect 333 120 338 132
rect 340 124 348 132
rect 340 122 343 124
rect 345 122 348 124
rect 340 120 348 122
rect 350 120 355 132
rect 357 130 364 132
rect 357 128 360 130
rect 362 128 364 130
rect 387 130 389 132
rect 391 130 394 132
rect 387 128 394 130
rect 357 126 364 128
rect 357 120 363 126
rect 299 117 306 119
rect 299 112 304 117
rect 359 118 363 120
rect 389 120 394 128
rect 396 120 401 140
rect 403 138 412 140
rect 618 139 627 141
rect 403 136 408 138
rect 410 136 412 138
rect 403 131 412 136
rect 618 137 621 139
rect 623 137 627 139
rect 403 129 408 131
rect 410 129 412 131
rect 403 126 412 129
rect 425 131 432 133
rect 425 129 427 131
rect 429 129 432 131
rect 425 127 432 129
rect 403 120 411 126
rect 359 112 365 118
rect 367 116 374 118
rect 367 114 370 116
rect 372 114 374 116
rect 367 112 374 114
rect 426 121 432 127
rect 434 121 439 133
rect 441 125 449 133
rect 441 123 444 125
rect 446 123 449 125
rect 441 121 449 123
rect 451 121 456 133
rect 458 131 466 133
rect 458 129 461 131
rect 463 129 466 131
rect 458 121 466 129
rect 468 127 473 133
rect 481 127 486 133
rect 468 125 475 127
rect 468 123 471 125
rect 473 123 475 125
rect 468 121 475 123
rect 479 125 486 127
rect 479 123 481 125
rect 483 123 486 125
rect 479 121 486 123
rect 488 131 496 133
rect 488 129 491 131
rect 493 129 496 131
rect 488 121 496 129
rect 498 121 503 133
rect 505 125 513 133
rect 505 123 508 125
rect 510 123 513 125
rect 505 121 513 123
rect 515 121 520 133
rect 522 131 529 133
rect 522 129 525 131
rect 527 129 529 131
rect 522 127 529 129
rect 522 121 528 127
rect 545 127 550 133
rect 426 119 430 121
rect 415 117 422 119
rect 415 115 417 117
rect 419 115 422 117
rect 415 113 422 115
rect 424 113 430 119
rect 524 119 528 121
rect 543 125 550 127
rect 543 123 545 125
rect 547 123 550 125
rect 543 121 550 123
rect 552 131 560 133
rect 552 129 555 131
rect 557 129 560 131
rect 552 121 560 129
rect 562 121 567 133
rect 569 125 577 133
rect 569 123 572 125
rect 574 123 577 125
rect 569 121 577 123
rect 579 121 584 133
rect 586 131 593 133
rect 618 132 627 137
rect 586 129 589 131
rect 591 129 593 131
rect 586 127 593 129
rect 607 130 614 132
rect 607 128 609 130
rect 611 128 614 130
rect 586 121 592 127
rect 607 126 614 128
rect 524 113 530 119
rect 532 117 539 119
rect 532 115 535 117
rect 537 115 539 117
rect 532 113 539 115
rect 588 119 592 121
rect 609 120 614 126
rect 616 123 627 132
rect 629 123 634 141
rect 636 134 641 141
rect 636 132 643 134
rect 636 130 639 132
rect 641 130 643 132
rect 636 128 643 130
rect 636 123 641 128
rect 616 120 624 123
rect 588 113 594 119
rect 596 117 603 119
rect 596 115 599 117
rect 601 115 603 117
rect 596 113 603 115
rect 650 119 655 125
rect 648 117 655 119
rect 648 115 650 117
rect 652 115 655 117
rect 648 113 655 115
rect 657 123 663 125
rect 657 117 665 123
rect 657 115 660 117
rect 662 115 665 117
rect 657 113 665 115
rect 667 117 675 123
rect 667 115 670 117
rect 672 115 675 117
rect 667 113 675 115
rect 677 121 684 123
rect 677 119 680 121
rect 682 119 684 121
rect 677 113 684 119
rect 4 27 11 33
rect 4 25 6 27
rect 8 25 11 27
rect 4 23 11 25
rect 13 31 21 33
rect 13 29 16 31
rect 18 29 21 31
rect 13 23 21 29
rect 23 31 31 33
rect 23 29 26 31
rect 28 29 31 31
rect 23 23 31 29
rect 25 21 31 23
rect 33 31 40 33
rect 33 29 36 31
rect 38 29 40 31
rect 33 27 40 29
rect 33 21 38 27
rect 85 31 92 33
rect 85 29 87 31
rect 89 29 92 31
rect 85 27 92 29
rect 94 27 100 33
rect 64 23 72 26
rect 47 18 52 23
rect 45 16 52 18
rect 45 14 47 16
rect 49 14 52 16
rect 45 12 52 14
rect 47 5 52 12
rect 54 5 59 23
rect 61 14 72 23
rect 74 20 79 26
rect 96 25 100 27
rect 149 31 156 33
rect 149 29 151 31
rect 153 29 156 31
rect 149 27 156 29
rect 158 27 164 33
rect 74 18 81 20
rect 96 19 102 25
rect 74 16 77 18
rect 79 16 81 18
rect 74 14 81 16
rect 95 17 102 19
rect 95 15 97 17
rect 99 15 102 17
rect 61 9 70 14
rect 95 13 102 15
rect 104 13 109 25
rect 111 23 119 25
rect 111 21 114 23
rect 116 21 119 23
rect 111 13 119 21
rect 121 13 126 25
rect 128 17 136 25
rect 128 15 131 17
rect 133 15 136 17
rect 128 13 136 15
rect 138 23 145 25
rect 138 21 141 23
rect 143 21 145 23
rect 138 19 145 21
rect 160 25 164 27
rect 258 27 264 33
rect 266 31 273 33
rect 266 29 269 31
rect 271 29 273 31
rect 266 27 273 29
rect 258 25 262 27
rect 138 13 143 19
rect 160 19 166 25
rect 159 17 166 19
rect 159 15 161 17
rect 163 15 166 17
rect 159 13 166 15
rect 168 13 173 25
rect 175 23 183 25
rect 175 21 178 23
rect 180 21 183 23
rect 175 13 183 21
rect 185 13 190 25
rect 192 17 200 25
rect 192 15 195 17
rect 197 15 200 17
rect 192 13 200 15
rect 202 23 209 25
rect 202 21 205 23
rect 207 21 209 23
rect 202 19 209 21
rect 213 23 220 25
rect 213 21 215 23
rect 217 21 220 23
rect 213 19 220 21
rect 202 13 207 19
rect 215 13 220 19
rect 222 17 230 25
rect 222 15 225 17
rect 227 15 230 17
rect 222 13 230 15
rect 232 13 237 25
rect 239 23 247 25
rect 239 21 242 23
rect 244 21 247 23
rect 239 13 247 21
rect 249 13 254 25
rect 256 19 262 25
rect 314 32 321 34
rect 314 30 316 32
rect 318 30 321 32
rect 314 28 321 30
rect 323 28 329 34
rect 277 20 285 26
rect 256 17 263 19
rect 256 15 259 17
rect 261 15 263 17
rect 256 13 263 15
rect 276 17 285 20
rect 276 15 278 17
rect 280 15 285 17
rect 61 7 65 9
rect 67 7 70 9
rect 276 10 285 15
rect 276 8 278 10
rect 280 8 285 10
rect 61 5 70 7
rect 276 6 285 8
rect 287 6 292 26
rect 294 18 299 26
rect 325 26 329 28
rect 384 29 389 34
rect 382 27 389 29
rect 325 20 331 26
rect 324 18 331 20
rect 294 16 301 18
rect 294 14 297 16
rect 299 14 301 16
rect 324 16 326 18
rect 328 16 331 18
rect 324 14 331 16
rect 333 14 338 26
rect 340 24 348 26
rect 340 22 343 24
rect 345 22 348 24
rect 340 14 348 22
rect 350 14 355 26
rect 357 18 365 26
rect 357 16 360 18
rect 362 16 365 18
rect 357 14 365 16
rect 367 24 374 26
rect 367 22 370 24
rect 372 22 374 24
rect 367 20 374 22
rect 382 25 384 27
rect 386 25 389 27
rect 382 20 389 25
rect 367 14 372 20
rect 382 18 384 20
rect 386 18 389 20
rect 382 16 389 18
rect 391 27 399 34
rect 423 32 430 34
rect 423 30 425 32
rect 427 30 430 32
rect 391 16 402 27
rect 294 12 301 14
rect 294 6 299 12
rect 393 10 402 16
rect 393 8 395 10
rect 397 8 402 10
rect 393 6 402 8
rect 404 6 409 27
rect 411 19 416 27
rect 423 25 430 30
rect 423 23 425 25
rect 427 23 430 25
rect 423 21 430 23
rect 411 17 418 19
rect 411 15 414 17
rect 416 15 418 17
rect 411 13 418 15
rect 411 6 416 13
rect 425 6 430 21
rect 432 17 440 34
rect 432 15 435 17
rect 437 15 440 17
rect 432 10 440 15
rect 432 8 435 10
rect 437 8 440 10
rect 432 6 440 8
rect 442 25 450 34
rect 442 23 445 25
rect 447 23 450 25
rect 442 18 450 23
rect 442 16 445 18
rect 447 16 450 18
rect 442 6 450 16
rect 452 17 468 34
rect 452 15 457 17
rect 459 15 468 17
rect 452 10 468 15
rect 452 8 457 10
rect 459 9 468 10
rect 470 9 475 34
rect 477 31 482 34
rect 512 32 519 34
rect 477 29 485 31
rect 477 27 480 29
rect 482 27 485 29
rect 477 18 485 27
rect 487 18 498 31
rect 477 9 482 18
rect 489 10 498 18
rect 459 8 466 9
rect 452 6 466 8
rect 489 8 492 10
rect 494 8 498 10
rect 489 6 498 8
rect 500 29 507 31
rect 500 27 503 29
rect 505 27 507 29
rect 500 22 507 27
rect 500 20 503 22
rect 505 20 507 22
rect 512 30 514 32
rect 516 30 519 32
rect 512 25 519 30
rect 512 23 514 25
rect 516 23 519 25
rect 512 21 519 23
rect 500 18 507 20
rect 500 6 505 18
rect 514 6 519 21
rect 521 17 529 34
rect 521 15 524 17
rect 526 15 529 17
rect 521 10 529 15
rect 521 8 524 10
rect 526 8 529 10
rect 521 6 529 8
rect 531 25 539 34
rect 531 23 534 25
rect 536 23 539 25
rect 531 18 539 23
rect 531 16 534 18
rect 536 16 539 18
rect 531 6 539 16
rect 541 17 557 34
rect 541 15 546 17
rect 548 15 557 17
rect 541 10 557 15
rect 541 8 546 10
rect 548 9 557 10
rect 559 9 564 34
rect 566 31 571 34
rect 600 32 607 34
rect 566 29 574 31
rect 566 27 569 29
rect 571 27 574 29
rect 566 18 574 27
rect 576 18 587 31
rect 566 9 571 18
rect 578 10 587 18
rect 548 8 555 9
rect 541 6 555 8
rect 578 8 581 10
rect 583 8 587 10
rect 578 6 587 8
rect 589 29 596 31
rect 589 27 592 29
rect 594 27 596 29
rect 600 30 602 32
rect 604 30 607 32
rect 600 28 607 30
rect 589 22 596 27
rect 602 26 607 28
rect 609 26 615 34
rect 589 20 592 22
rect 594 20 596 22
rect 589 18 596 20
rect 611 22 615 26
rect 664 32 671 34
rect 664 30 666 32
rect 668 30 671 32
rect 664 25 671 30
rect 646 22 651 24
rect 589 6 594 18
rect 611 18 617 22
rect 610 10 617 18
rect 610 8 612 10
rect 614 8 617 10
rect 610 6 617 8
rect 619 6 624 22
rect 626 20 634 22
rect 626 18 629 20
rect 631 18 634 20
rect 626 6 634 18
rect 636 6 641 22
rect 643 10 651 22
rect 643 8 646 10
rect 648 8 651 10
rect 643 6 651 8
rect 653 19 658 24
rect 664 23 666 25
rect 668 23 671 25
rect 664 21 671 23
rect 653 17 660 19
rect 653 15 656 17
rect 658 15 660 17
rect 666 16 671 21
rect 673 17 682 34
rect 673 16 677 17
rect 653 13 660 15
rect 653 6 658 13
rect 675 15 677 16
rect 679 15 682 17
rect 675 13 682 15
<< alu1 >>
rect -16 290 688 293
rect -18 289 688 290
rect -18 288 418 289
rect -18 286 7 288
rect 9 286 19 288
rect 21 286 301 288
rect 303 286 369 288
rect 371 287 418 288
rect 420 287 534 289
rect 536 287 598 289
rect 600 287 610 289
rect 612 287 651 289
rect 653 287 665 289
rect 667 287 679 289
rect 681 287 688 289
rect 371 286 688 287
rect -18 285 412 286
rect -18 150 -11 285
rect 28 278 41 279
rect 28 276 30 278
rect 32 276 41 278
rect 28 275 41 276
rect 12 270 24 272
rect 12 268 20 270
rect 22 268 24 270
rect 12 266 24 268
rect 20 263 24 266
rect 22 261 24 263
rect 4 254 16 256
rect 4 252 6 254
rect 8 252 13 254
rect 15 252 16 254
rect 4 250 16 252
rect 12 242 16 250
rect 20 249 24 261
rect 20 247 21 249
rect 23 247 24 249
rect 20 245 24 247
rect 22 243 24 245
rect 20 234 24 243
rect 28 254 32 275
rect 83 274 88 280
rect 83 272 84 274
rect 86 272 88 274
rect 28 252 29 254
rect 31 252 32 254
rect 28 242 32 252
rect 83 271 88 272
rect 75 267 88 271
rect 92 275 105 279
rect 181 275 194 279
rect 302 279 306 280
rect 293 275 306 279
rect 92 273 97 275
rect 92 271 94 273
rect 96 271 97 273
rect 181 273 186 275
rect 92 266 97 271
rect 92 264 94 266
rect 96 264 97 266
rect 44 262 56 264
rect 44 260 49 262
rect 51 260 56 262
rect 44 259 56 260
rect 46 258 56 259
rect 46 257 48 258
rect 44 250 48 257
rect 68 254 74 256
rect 68 252 71 254
rect 73 252 74 254
rect 68 247 74 252
rect 68 246 81 247
rect 68 244 69 246
rect 71 244 81 246
rect 68 243 81 244
rect 28 240 33 242
rect 28 238 30 240
rect 32 238 33 240
rect 28 236 33 238
rect 28 234 32 236
rect 92 262 97 264
rect 92 242 96 262
rect 123 262 161 263
rect 123 260 152 262
rect 154 260 161 262
rect 123 259 161 260
rect 123 256 128 259
rect 120 254 128 256
rect 120 252 121 254
rect 123 252 128 254
rect 120 250 128 252
rect 138 254 153 255
rect 138 252 140 254
rect 142 252 147 254
rect 149 252 153 254
rect 138 251 153 252
rect 92 240 93 242
rect 95 240 96 242
rect 92 238 97 240
rect 140 245 144 251
rect 171 270 177 272
rect 171 268 172 270
rect 174 268 177 270
rect 171 263 177 268
rect 171 261 172 263
rect 174 261 177 263
rect 171 259 177 261
rect 140 243 141 245
rect 143 243 144 245
rect 140 242 144 243
rect 173 245 177 259
rect 173 243 174 245
rect 176 243 177 245
rect 173 239 177 243
rect 92 236 94 238
rect 96 236 97 238
rect 92 234 97 236
rect 155 238 177 239
rect 155 236 172 238
rect 174 236 177 238
rect 155 235 177 236
rect 181 271 183 273
rect 185 271 186 273
rect 181 266 186 271
rect 181 264 183 266
rect 185 264 186 266
rect 181 262 186 264
rect 181 260 182 262
rect 184 260 185 262
rect 181 240 185 260
rect 212 259 250 263
rect 212 256 217 259
rect 209 254 217 256
rect 209 252 210 254
rect 212 252 214 254
rect 216 252 217 254
rect 209 250 217 252
rect 227 254 242 255
rect 227 252 229 254
rect 231 252 236 254
rect 238 252 242 254
rect 227 251 242 252
rect 181 238 186 240
rect 229 242 233 251
rect 260 270 266 272
rect 260 268 261 270
rect 263 269 266 270
rect 270 269 274 272
rect 263 268 274 269
rect 260 265 274 268
rect 260 263 266 265
rect 260 261 261 263
rect 263 261 266 263
rect 260 259 266 261
rect 270 263 274 265
rect 270 261 291 263
rect 270 259 275 261
rect 277 259 291 261
rect 262 239 266 259
rect 270 254 291 255
rect 270 252 285 254
rect 287 252 291 254
rect 270 251 291 252
rect 304 273 306 275
rect 369 278 374 280
rect 369 276 370 278
rect 372 276 374 278
rect 302 268 306 273
rect 369 272 374 276
rect 304 266 306 268
rect 270 245 274 251
rect 302 256 306 266
rect 302 254 303 256
rect 305 254 306 256
rect 302 247 306 254
rect 270 243 271 245
rect 273 243 274 245
rect 270 242 274 243
rect 301 245 306 247
rect 301 243 302 245
rect 304 243 306 245
rect 301 241 306 243
rect 314 271 320 272
rect 369 271 370 272
rect 314 269 316 271
rect 318 269 327 271
rect 314 267 327 269
rect 361 270 370 271
rect 372 270 374 272
rect 361 267 374 270
rect 384 279 393 280
rect 384 277 389 279
rect 391 277 393 279
rect 384 276 393 277
rect 181 236 183 238
rect 185 236 186 238
rect 181 234 186 236
rect 244 238 266 239
rect 244 236 261 238
rect 263 236 266 238
rect 244 235 266 236
rect 314 238 318 267
rect 337 257 343 263
rect 328 256 343 257
rect 328 254 330 256
rect 332 254 339 256
rect 341 254 343 256
rect 328 251 343 254
rect 354 254 360 256
rect 354 252 357 254
rect 359 252 360 254
rect 354 248 360 252
rect 354 245 366 248
rect 354 243 360 245
rect 362 243 366 245
rect 354 242 366 243
rect 314 237 320 238
rect 314 235 316 237
rect 318 235 320 237
rect 314 234 320 235
rect 384 259 388 276
rect 415 278 420 280
rect 415 276 416 278
rect 418 276 420 278
rect 415 273 420 276
rect 534 277 539 281
rect 534 275 536 277
rect 538 275 539 277
rect 603 285 607 286
rect 598 278 603 281
rect 598 276 600 278
rect 602 276 603 278
rect 534 273 539 275
rect 598 273 603 276
rect 400 271 404 272
rect 400 269 401 271
rect 403 269 404 271
rect 400 267 404 269
rect 415 271 417 273
rect 419 272 420 273
rect 469 272 475 273
rect 419 271 428 272
rect 415 268 428 271
rect 462 270 471 272
rect 473 270 475 272
rect 462 268 475 270
rect 384 257 385 259
rect 387 257 388 259
rect 392 263 404 267
rect 408 263 412 264
rect 392 262 396 263
rect 392 260 393 262
rect 395 260 396 262
rect 392 258 396 260
rect 408 261 409 263
rect 411 261 412 263
rect 384 254 388 257
rect 408 256 412 261
rect 384 250 396 254
rect 400 253 412 256
rect 400 251 403 253
rect 405 251 412 253
rect 400 250 412 251
rect 392 245 396 250
rect 392 244 401 245
rect 392 242 397 244
rect 399 242 401 244
rect 392 241 401 242
rect 429 255 435 257
rect 429 253 430 255
rect 432 253 435 255
rect 429 249 435 253
rect 423 247 435 249
rect 423 245 429 247
rect 431 245 435 247
rect 423 243 435 245
rect 446 258 452 264
rect 446 257 461 258
rect 446 256 457 257
rect 446 254 452 256
rect 454 255 457 256
rect 459 255 461 257
rect 454 254 461 255
rect 446 252 461 254
rect 471 256 475 268
rect 471 254 472 256
rect 474 254 475 256
rect 471 239 475 254
rect 469 238 475 239
rect 469 236 471 238
rect 473 236 475 238
rect 469 235 475 236
rect 479 272 485 273
rect 534 272 535 273
rect 479 270 481 272
rect 483 270 492 272
rect 479 268 492 270
rect 526 271 535 272
rect 537 271 539 273
rect 526 268 539 271
rect 543 272 549 273
rect 598 272 599 273
rect 543 270 545 272
rect 547 270 556 272
rect 543 268 556 270
rect 590 271 599 272
rect 601 271 603 273
rect 590 268 603 271
rect 607 277 620 280
rect 607 275 609 277
rect 611 276 620 277
rect 479 239 483 268
rect 502 258 508 264
rect 493 257 508 258
rect 493 255 495 257
rect 497 256 508 257
rect 497 255 500 256
rect 493 254 500 255
rect 502 254 508 256
rect 493 252 508 254
rect 519 255 525 257
rect 519 253 522 255
rect 524 253 525 255
rect 519 249 525 253
rect 519 247 531 249
rect 519 245 524 247
rect 526 245 531 247
rect 519 243 531 245
rect 479 238 485 239
rect 479 236 481 238
rect 483 236 485 238
rect 479 235 485 236
rect 543 247 547 268
rect 543 245 544 247
rect 546 245 547 247
rect 543 239 547 245
rect 566 259 572 264
rect 566 258 569 259
rect 557 257 569 258
rect 571 257 572 259
rect 557 255 559 257
rect 561 255 572 257
rect 557 252 572 255
rect 583 255 589 257
rect 583 253 586 255
rect 588 253 589 255
rect 583 249 589 253
rect 583 246 595 249
rect 583 244 592 246
rect 594 244 595 246
rect 583 243 595 244
rect 543 238 549 239
rect 543 236 545 238
rect 547 236 549 238
rect 543 235 549 236
rect 607 259 611 275
rect 607 257 608 259
rect 610 257 611 259
rect 607 243 611 257
rect 631 272 635 273
rect 631 270 632 272
rect 634 270 635 272
rect 631 264 635 270
rect 622 263 635 264
rect 622 261 626 263
rect 628 261 635 263
rect 622 260 635 261
rect 639 256 643 265
rect 630 255 643 256
rect 630 253 636 255
rect 638 253 640 255
rect 642 253 643 255
rect 630 252 643 253
rect 639 251 643 252
rect 648 264 652 273
rect 648 262 650 264
rect 607 241 612 243
rect 607 239 609 241
rect 611 239 612 241
rect 607 235 612 239
rect 648 246 652 262
rect 663 279 691 281
rect 663 277 667 279
rect 669 277 691 279
rect 663 275 676 277
rect 663 272 669 275
rect 663 270 665 272
rect 667 270 669 272
rect 663 268 669 270
rect 680 255 684 257
rect 680 253 681 255
rect 683 253 684 255
rect 648 244 649 246
rect 651 244 652 246
rect 648 241 652 244
rect 648 239 650 241
rect 652 239 660 241
rect 648 235 660 239
rect 680 251 684 253
rect 680 248 693 251
rect 671 247 693 248
rect 671 245 676 247
rect 678 245 684 247
rect 671 243 684 245
rect 383 229 688 230
rect 0 228 610 229
rect 0 226 7 228
rect 9 226 19 228
rect 21 226 301 228
rect 303 226 387 228
rect 389 226 407 228
rect 409 227 610 228
rect 612 227 638 229
rect 640 227 651 229
rect 653 227 661 229
rect 663 227 688 229
rect 409 226 688 227
rect 0 214 708 226
rect 0 213 279 214
rect 0 211 25 213
rect 27 211 35 213
rect 37 211 48 213
rect 50 211 76 213
rect 78 212 279 213
rect 281 212 299 214
rect 301 212 385 214
rect 387 212 667 214
rect 669 212 679 214
rect 681 212 688 214
rect 78 211 688 212
rect 0 210 306 211
rect 4 195 17 197
rect 4 193 10 195
rect 12 193 17 195
rect 4 192 17 193
rect 4 187 8 192
rect 28 201 40 205
rect 28 199 36 201
rect 38 199 40 201
rect 36 196 40 199
rect 36 194 37 196
rect 39 194 40 196
rect 4 185 5 187
rect 7 185 8 187
rect 4 183 8 185
rect 19 170 25 172
rect 19 168 21 170
rect 23 168 25 170
rect 19 165 25 168
rect 12 163 25 165
rect 12 161 19 163
rect 21 161 25 163
rect 12 159 25 161
rect 36 178 40 194
rect 76 201 81 205
rect 76 199 77 201
rect 79 199 81 201
rect 76 197 81 199
rect 38 176 40 178
rect 36 167 40 176
rect 45 188 49 189
rect 45 187 58 188
rect 45 185 46 187
rect 48 185 50 187
rect 52 185 58 187
rect 45 184 58 185
rect 45 175 49 184
rect 53 179 66 180
rect 53 177 60 179
rect 62 177 66 179
rect 53 176 66 177
rect 53 170 57 176
rect 53 168 54 170
rect 56 168 57 170
rect 53 167 57 168
rect 77 183 81 197
rect 77 181 78 183
rect 80 181 81 183
rect 77 165 81 181
rect 139 204 145 205
rect 139 202 141 204
rect 143 202 145 204
rect 139 201 145 202
rect 93 196 105 197
rect 93 194 94 196
rect 96 194 105 196
rect 93 191 105 194
rect 99 187 105 191
rect 99 185 100 187
rect 102 185 105 187
rect 99 183 105 185
rect 116 185 131 188
rect 116 183 127 185
rect 129 183 131 185
rect 116 181 117 183
rect 119 182 131 183
rect 119 181 122 182
rect 116 176 122 181
rect 141 195 145 201
rect 141 193 142 195
rect 144 193 145 195
rect 141 172 145 193
rect 203 204 209 205
rect 203 202 205 204
rect 207 202 209 204
rect 203 201 209 202
rect 157 195 169 197
rect 157 193 162 195
rect 164 193 169 195
rect 157 191 169 193
rect 163 187 169 191
rect 163 185 164 187
rect 166 185 169 187
rect 163 183 169 185
rect 180 186 195 188
rect 180 184 186 186
rect 188 185 195 186
rect 188 184 191 185
rect 180 183 191 184
rect 193 183 195 185
rect 180 182 195 183
rect 180 176 186 182
rect 205 172 209 201
rect 68 163 77 164
rect 79 163 81 165
rect 68 160 81 163
rect 85 169 98 172
rect 85 167 87 169
rect 89 168 98 169
rect 132 170 145 172
rect 132 168 141 170
rect 143 168 145 170
rect 89 167 90 168
rect 139 167 145 168
rect 149 169 162 172
rect 149 167 151 169
rect 153 168 162 169
rect 196 170 209 172
rect 196 168 205 170
rect 207 168 209 170
rect 153 167 154 168
rect 203 167 209 168
rect 213 204 219 205
rect 213 202 215 204
rect 217 202 219 204
rect 213 201 219 202
rect 213 186 217 201
rect 213 184 214 186
rect 216 184 217 186
rect 213 172 217 184
rect 227 186 242 188
rect 227 185 234 186
rect 227 183 229 185
rect 231 184 234 185
rect 236 184 242 186
rect 231 183 242 184
rect 227 182 242 183
rect 236 176 242 182
rect 253 195 265 197
rect 253 193 257 195
rect 259 193 265 195
rect 253 191 265 193
rect 253 187 259 191
rect 253 185 256 187
rect 258 185 259 187
rect 253 183 259 185
rect 287 198 296 199
rect 287 196 289 198
rect 291 196 296 198
rect 287 195 296 196
rect 292 190 296 195
rect 276 189 288 190
rect 276 187 283 189
rect 285 187 288 189
rect 276 184 288 187
rect 292 186 304 190
rect 276 179 280 184
rect 300 183 304 186
rect 276 177 277 179
rect 279 177 280 179
rect 292 180 296 182
rect 292 178 293 180
rect 295 178 296 180
rect 292 177 296 178
rect 276 176 280 177
rect 284 173 296 177
rect 300 181 301 183
rect 303 181 304 183
rect 213 170 226 172
rect 213 168 215 170
rect 217 168 226 170
rect 260 169 273 172
rect 260 168 269 169
rect 213 167 219 168
rect 268 167 269 168
rect 271 167 273 169
rect 284 171 288 173
rect 284 169 285 171
rect 287 169 288 171
rect 284 168 288 169
rect 85 164 90 167
rect 149 165 154 167
rect 85 162 86 164
rect 88 162 90 164
rect 85 159 90 162
rect 81 154 85 155
rect 149 163 150 165
rect 152 163 154 165
rect 149 159 154 163
rect 268 164 273 167
rect 268 162 270 164
rect 272 162 273 164
rect 268 160 273 162
rect 300 164 304 181
rect 368 205 374 206
rect 368 203 370 205
rect 372 203 374 205
rect 368 202 374 203
rect 322 197 334 198
rect 322 195 326 197
rect 328 195 334 197
rect 322 192 334 195
rect 328 188 334 192
rect 328 186 329 188
rect 331 186 334 188
rect 328 184 334 186
rect 345 186 360 189
rect 345 184 347 186
rect 349 184 356 186
rect 358 184 360 186
rect 345 183 360 184
rect 345 177 351 183
rect 370 178 374 202
rect 422 204 444 205
rect 422 202 425 204
rect 427 202 444 204
rect 422 201 444 202
rect 502 204 507 206
rect 502 202 503 204
rect 505 202 507 204
rect 370 176 371 178
rect 373 176 374 178
rect 370 173 374 176
rect 295 163 304 164
rect 295 161 297 163
rect 299 161 304 163
rect 295 160 304 161
rect 314 170 327 173
rect 314 168 316 170
rect 318 169 327 170
rect 361 171 374 173
rect 361 169 370 171
rect 372 169 374 171
rect 318 168 319 169
rect 368 168 374 169
rect 382 197 387 199
rect 382 195 384 197
rect 386 195 387 197
rect 382 193 387 195
rect 414 197 418 198
rect 414 195 415 197
rect 417 195 418 197
rect 382 186 386 193
rect 382 184 383 186
rect 385 184 386 186
rect 382 174 386 184
rect 414 189 418 195
rect 382 172 384 174
rect 314 164 319 168
rect 382 167 386 172
rect 314 162 316 164
rect 318 162 319 164
rect 314 160 319 162
rect 382 165 384 167
rect 397 188 418 189
rect 397 186 401 188
rect 403 186 418 188
rect 397 185 418 186
rect 422 181 426 201
rect 397 179 411 181
rect 413 179 418 181
rect 397 177 418 179
rect 414 175 418 177
rect 422 179 428 181
rect 422 177 425 179
rect 427 177 428 179
rect 422 175 428 177
rect 414 172 428 175
rect 414 171 425 172
rect 414 168 418 171
rect 422 170 425 171
rect 427 170 428 172
rect 422 168 428 170
rect 455 189 459 198
rect 502 200 507 202
rect 446 188 461 189
rect 446 186 450 188
rect 452 186 457 188
rect 459 186 461 188
rect 446 185 461 186
rect 471 188 479 190
rect 471 186 472 188
rect 474 186 476 188
rect 478 186 479 188
rect 471 184 479 186
rect 471 181 476 184
rect 438 177 476 181
rect 503 180 507 200
rect 503 178 504 180
rect 506 178 507 180
rect 502 176 507 178
rect 502 174 503 176
rect 505 174 507 176
rect 502 169 507 174
rect 502 167 503 169
rect 505 167 507 169
rect 511 204 533 205
rect 511 202 514 204
rect 516 202 533 204
rect 511 201 533 202
rect 591 204 596 206
rect 591 202 592 204
rect 594 202 596 204
rect 511 197 515 201
rect 511 195 512 197
rect 514 195 515 197
rect 511 181 515 195
rect 544 197 548 198
rect 544 195 545 197
rect 547 195 548 197
rect 511 179 517 181
rect 511 177 514 179
rect 516 177 517 179
rect 511 172 517 177
rect 511 170 514 172
rect 516 170 517 172
rect 511 168 517 170
rect 544 189 548 195
rect 591 200 596 202
rect 592 198 593 200
rect 595 198 596 200
rect 535 188 550 189
rect 535 186 539 188
rect 541 186 546 188
rect 548 186 550 188
rect 535 185 550 186
rect 560 188 568 190
rect 560 186 565 188
rect 567 186 568 188
rect 560 184 568 186
rect 560 181 565 184
rect 527 180 565 181
rect 527 178 534 180
rect 536 178 565 180
rect 527 177 565 178
rect 592 178 596 198
rect 591 176 596 178
rect 656 204 660 206
rect 655 202 660 204
rect 655 200 656 202
rect 658 200 660 202
rect 655 198 660 200
rect 607 196 620 197
rect 607 194 617 196
rect 619 194 620 196
rect 607 193 620 194
rect 614 188 620 193
rect 614 186 615 188
rect 617 186 620 188
rect 614 184 620 186
rect 640 183 644 190
rect 640 182 642 183
rect 632 181 642 182
rect 632 180 644 181
rect 632 178 637 180
rect 639 178 644 180
rect 632 176 644 178
rect 591 174 592 176
rect 594 174 596 176
rect 591 169 596 174
rect 502 165 507 167
rect 591 167 592 169
rect 594 167 596 169
rect 591 165 596 167
rect 382 161 395 165
rect 382 160 386 161
rect 494 161 507 165
rect 583 161 596 165
rect 600 171 613 173
rect 600 169 602 171
rect 604 169 613 171
rect 600 168 605 169
rect 656 188 660 198
rect 656 186 657 188
rect 659 186 660 188
rect 600 166 602 168
rect 604 166 605 168
rect 600 160 605 166
rect 656 165 660 186
rect 664 197 668 206
rect 664 195 666 197
rect 664 193 668 195
rect 664 191 665 193
rect 667 191 668 193
rect 664 179 668 191
rect 672 190 676 198
rect 672 188 684 190
rect 672 186 673 188
rect 675 186 680 188
rect 682 186 684 188
rect 672 184 684 186
rect 664 177 666 179
rect 664 174 668 177
rect 664 172 676 174
rect 664 170 666 172
rect 668 170 676 172
rect 664 168 676 170
rect 647 164 660 165
rect 647 162 656 164
rect 658 162 660 164
rect 647 161 660 162
rect 276 154 688 155
rect 0 153 317 154
rect 0 151 7 153
rect 9 151 21 153
rect 23 151 35 153
rect 37 151 76 153
rect 78 151 88 153
rect 90 151 152 153
rect 154 151 268 153
rect 270 152 317 153
rect 319 152 385 154
rect 387 152 667 154
rect 669 152 679 154
rect 681 152 688 154
rect 270 151 688 152
rect 0 150 688 151
rect -18 142 688 150
rect -18 8 -11 142
rect 0 141 418 142
rect 0 139 7 141
rect 9 139 19 141
rect 21 139 301 141
rect 303 139 369 141
rect 371 140 418 141
rect 420 140 534 142
rect 536 140 598 142
rect 600 140 610 142
rect 612 140 651 142
rect 653 140 665 142
rect 667 140 679 142
rect 681 140 688 142
rect 371 139 688 140
rect 0 138 412 139
rect 28 131 41 132
rect 28 129 30 131
rect 32 129 41 131
rect 28 128 41 129
rect 12 123 24 125
rect 12 121 20 123
rect 22 121 24 123
rect 12 119 24 121
rect 20 116 24 119
rect 22 114 24 116
rect 4 107 16 109
rect 4 105 6 107
rect 8 105 13 107
rect 15 105 16 107
rect 4 103 16 105
rect 12 95 16 103
rect 20 102 24 114
rect 20 100 21 102
rect 23 100 24 102
rect 20 98 24 100
rect 22 96 24 98
rect 20 87 24 96
rect 28 107 32 128
rect 83 127 88 133
rect 83 125 84 127
rect 86 125 88 127
rect 28 105 29 107
rect 31 105 32 107
rect 28 95 32 105
rect 83 124 88 125
rect 75 120 88 124
rect 92 128 105 132
rect 181 128 194 132
rect 302 132 306 133
rect 293 128 306 132
rect 92 126 97 128
rect 92 124 94 126
rect 96 124 97 126
rect 181 126 186 128
rect 92 119 97 124
rect 92 117 94 119
rect 96 117 97 119
rect 44 115 56 117
rect 44 113 49 115
rect 51 113 56 115
rect 44 112 56 113
rect 46 111 56 112
rect 46 110 48 111
rect 44 103 48 110
rect 68 107 74 109
rect 68 105 71 107
rect 73 105 74 107
rect 68 100 74 105
rect 68 99 81 100
rect 68 97 69 99
rect 71 97 81 99
rect 68 96 81 97
rect 28 93 33 95
rect 28 91 30 93
rect 32 91 33 93
rect 28 89 33 91
rect 28 87 32 89
rect 92 115 97 117
rect 92 95 96 115
rect 123 115 161 116
rect 123 113 152 115
rect 154 113 161 115
rect 123 112 161 113
rect 123 109 128 112
rect 120 107 128 109
rect 120 105 121 107
rect 123 105 128 107
rect 120 103 128 105
rect 138 107 153 108
rect 138 105 140 107
rect 142 105 147 107
rect 149 105 153 107
rect 138 104 153 105
rect 92 93 93 95
rect 95 93 96 95
rect 92 91 97 93
rect 140 98 144 104
rect 171 123 177 125
rect 171 121 172 123
rect 174 121 177 123
rect 171 116 177 121
rect 171 114 172 116
rect 174 114 177 116
rect 171 112 177 114
rect 140 96 141 98
rect 143 96 144 98
rect 140 95 144 96
rect 173 98 177 112
rect 173 96 174 98
rect 176 96 177 98
rect 173 92 177 96
rect 92 89 94 91
rect 96 89 97 91
rect 92 87 97 89
rect 155 91 177 92
rect 155 89 172 91
rect 174 89 177 91
rect 155 88 177 89
rect 181 124 183 126
rect 185 124 186 126
rect 181 119 186 124
rect 181 117 183 119
rect 185 117 186 119
rect 181 115 186 117
rect 181 113 182 115
rect 184 113 185 115
rect 181 93 185 113
rect 212 112 250 116
rect 212 109 217 112
rect 209 107 217 109
rect 209 105 210 107
rect 212 105 214 107
rect 216 105 217 107
rect 209 103 217 105
rect 227 107 242 108
rect 227 105 229 107
rect 231 105 236 107
rect 238 105 242 107
rect 227 104 242 105
rect 181 91 186 93
rect 229 95 233 104
rect 260 123 266 125
rect 260 121 261 123
rect 263 122 266 123
rect 270 122 274 125
rect 263 121 274 122
rect 260 118 274 121
rect 260 116 266 118
rect 260 114 261 116
rect 263 114 266 116
rect 260 112 266 114
rect 270 116 274 118
rect 270 114 291 116
rect 270 112 275 114
rect 277 112 291 114
rect 262 92 266 112
rect 270 107 291 108
rect 270 105 285 107
rect 287 105 291 107
rect 270 104 291 105
rect 304 126 306 128
rect 369 131 374 133
rect 369 129 370 131
rect 372 129 374 131
rect 302 121 306 126
rect 369 125 374 129
rect 304 119 306 121
rect 270 98 274 104
rect 302 109 306 119
rect 302 107 303 109
rect 305 107 306 109
rect 302 100 306 107
rect 270 96 271 98
rect 273 96 274 98
rect 270 95 274 96
rect 301 98 306 100
rect 301 96 302 98
rect 304 96 306 98
rect 301 94 306 96
rect 314 124 320 125
rect 369 124 370 125
rect 314 122 316 124
rect 318 122 327 124
rect 314 120 327 122
rect 361 123 370 124
rect 372 123 374 125
rect 361 120 374 123
rect 384 132 393 133
rect 384 130 389 132
rect 391 130 393 132
rect 384 129 393 130
rect 181 89 183 91
rect 185 89 186 91
rect 181 87 186 89
rect 244 91 266 92
rect 244 89 261 91
rect 263 89 266 91
rect 244 88 266 89
rect 314 91 318 120
rect 337 110 343 116
rect 328 109 343 110
rect 328 107 330 109
rect 332 107 339 109
rect 341 107 343 109
rect 328 104 343 107
rect 354 107 360 109
rect 354 105 357 107
rect 359 105 360 107
rect 354 101 360 105
rect 354 98 366 101
rect 354 96 360 98
rect 362 96 366 98
rect 354 95 366 96
rect 314 90 320 91
rect 314 88 316 90
rect 318 88 320 90
rect 314 87 320 88
rect 384 112 388 129
rect 415 131 420 133
rect 415 129 416 131
rect 418 129 420 131
rect 415 126 420 129
rect 534 130 539 134
rect 534 128 536 130
rect 538 128 539 130
rect 603 138 607 139
rect 598 131 603 134
rect 598 129 600 131
rect 602 129 603 131
rect 534 126 539 128
rect 598 126 603 129
rect 400 124 404 125
rect 400 122 401 124
rect 403 122 404 124
rect 400 120 404 122
rect 415 124 417 126
rect 419 125 420 126
rect 469 125 475 126
rect 419 124 428 125
rect 415 121 428 124
rect 462 123 471 125
rect 473 123 475 125
rect 462 121 475 123
rect 384 110 385 112
rect 387 110 388 112
rect 392 116 404 120
rect 408 116 412 117
rect 392 115 396 116
rect 392 113 393 115
rect 395 113 396 115
rect 392 111 396 113
rect 408 114 409 116
rect 411 114 412 116
rect 384 107 388 110
rect 408 109 412 114
rect 384 103 396 107
rect 400 106 412 109
rect 400 104 403 106
rect 405 104 412 106
rect 400 103 412 104
rect 392 98 396 103
rect 392 97 401 98
rect 392 95 397 97
rect 399 95 401 97
rect 392 94 401 95
rect 429 108 435 110
rect 429 106 430 108
rect 432 106 435 108
rect 429 102 435 106
rect 423 100 435 102
rect 423 98 429 100
rect 431 98 435 100
rect 423 96 435 98
rect 446 111 452 117
rect 446 110 461 111
rect 446 109 457 110
rect 446 107 452 109
rect 454 108 457 109
rect 459 108 461 110
rect 454 107 461 108
rect 446 105 461 107
rect 471 109 475 121
rect 471 107 472 109
rect 474 107 475 109
rect 471 92 475 107
rect 469 91 475 92
rect 469 89 471 91
rect 473 89 475 91
rect 469 88 475 89
rect 479 125 485 126
rect 534 125 535 126
rect 479 123 481 125
rect 483 123 492 125
rect 479 121 492 123
rect 526 124 535 125
rect 537 124 539 126
rect 526 121 539 124
rect 543 125 549 126
rect 598 125 599 126
rect 543 123 545 125
rect 547 123 556 125
rect 543 121 556 123
rect 590 124 599 125
rect 601 124 603 126
rect 590 121 603 124
rect 607 130 620 133
rect 607 128 609 130
rect 611 129 620 130
rect 479 92 483 121
rect 502 111 508 117
rect 493 110 508 111
rect 493 108 495 110
rect 497 109 508 110
rect 497 108 500 109
rect 493 107 500 108
rect 502 107 508 109
rect 493 105 508 107
rect 519 108 525 110
rect 519 106 522 108
rect 524 106 525 108
rect 519 102 525 106
rect 519 100 531 102
rect 519 98 524 100
rect 526 98 531 100
rect 519 96 531 98
rect 479 91 485 92
rect 479 89 481 91
rect 483 89 485 91
rect 479 88 485 89
rect 543 100 547 121
rect 543 98 544 100
rect 546 98 547 100
rect 543 92 547 98
rect 566 112 572 117
rect 566 111 569 112
rect 557 110 569 111
rect 571 110 572 112
rect 557 108 559 110
rect 561 108 572 110
rect 557 105 572 108
rect 583 108 589 110
rect 583 106 586 108
rect 588 106 589 108
rect 583 102 589 106
rect 583 99 595 102
rect 583 97 592 99
rect 594 97 595 99
rect 583 96 595 97
rect 543 91 549 92
rect 543 89 545 91
rect 547 89 549 91
rect 543 88 549 89
rect 607 112 611 128
rect 607 110 608 112
rect 610 110 611 112
rect 607 96 611 110
rect 631 125 635 126
rect 631 123 632 125
rect 634 123 635 125
rect 631 117 635 123
rect 622 116 635 117
rect 622 114 626 116
rect 628 114 635 116
rect 622 113 635 114
rect 639 109 643 118
rect 630 108 643 109
rect 630 106 636 108
rect 638 106 640 108
rect 642 106 643 108
rect 630 105 643 106
rect 639 104 643 105
rect 648 117 652 126
rect 648 115 650 117
rect 607 94 612 96
rect 607 92 609 94
rect 611 92 612 94
rect 607 88 612 92
rect 648 99 652 115
rect 663 132 676 134
rect 663 130 667 132
rect 669 130 676 132
rect 663 128 676 130
rect 663 125 669 128
rect 663 123 665 125
rect 667 123 669 125
rect 663 121 669 123
rect 680 108 684 110
rect 680 106 681 108
rect 683 106 684 108
rect 648 97 649 99
rect 651 97 652 99
rect 648 94 652 97
rect 648 92 650 94
rect 652 92 660 94
rect 648 88 660 92
rect 680 101 684 106
rect 671 100 684 101
rect 671 98 676 100
rect 678 98 684 100
rect 671 96 684 98
rect 382 82 688 83
rect 0 81 610 82
rect 0 79 7 81
rect 9 79 19 81
rect 21 79 301 81
rect 303 79 387 81
rect 389 79 407 81
rect 409 80 610 81
rect 612 80 638 82
rect 640 80 651 82
rect 653 80 661 82
rect 663 81 688 82
rect 700 81 708 214
rect 663 80 708 81
rect 409 79 708 80
rect 0 69 708 79
rect 0 67 688 69
rect 0 66 279 67
rect 0 64 25 66
rect 27 64 35 66
rect 37 64 48 66
rect 50 64 76 66
rect 78 65 279 66
rect 281 65 299 67
rect 301 65 385 67
rect 387 65 667 67
rect 669 65 679 67
rect 681 65 688 67
rect 78 64 688 65
rect 0 63 305 64
rect 4 48 17 50
rect 4 46 10 48
rect 12 46 17 48
rect 4 45 17 46
rect 4 40 8 45
rect 28 54 40 58
rect 28 52 36 54
rect 38 52 40 54
rect 36 49 40 52
rect 36 47 37 49
rect 39 47 40 49
rect 4 38 5 40
rect 7 38 8 40
rect 4 36 8 38
rect -18 7 0 8
rect 19 23 25 25
rect 19 21 21 23
rect 23 21 25 23
rect 19 18 25 21
rect 12 16 25 18
rect 12 14 19 16
rect 21 14 25 16
rect 12 12 25 14
rect 36 31 40 47
rect 76 54 81 58
rect 76 52 77 54
rect 79 52 81 54
rect 76 50 81 52
rect 38 29 40 31
rect 36 20 40 29
rect 45 41 49 42
rect 45 40 58 41
rect 45 38 46 40
rect 48 38 50 40
rect 52 38 58 40
rect 45 37 58 38
rect 45 28 49 37
rect 53 32 66 33
rect 53 30 60 32
rect 62 30 66 32
rect 53 29 66 30
rect 53 23 57 29
rect 53 21 54 23
rect 56 21 57 23
rect 53 20 57 21
rect 77 36 81 50
rect 77 34 78 36
rect 80 34 81 36
rect 77 18 81 34
rect 139 57 145 58
rect 139 55 141 57
rect 143 55 145 57
rect 139 54 145 55
rect 93 49 105 50
rect 93 47 94 49
rect 96 47 105 49
rect 93 44 105 47
rect 99 40 105 44
rect 99 38 100 40
rect 102 38 105 40
rect 99 36 105 38
rect 116 38 131 41
rect 116 36 127 38
rect 129 36 131 38
rect 116 34 117 36
rect 119 35 131 36
rect 119 34 122 35
rect 116 29 122 34
rect 141 48 145 54
rect 141 46 142 48
rect 144 46 145 48
rect 141 25 145 46
rect 203 57 209 58
rect 203 55 205 57
rect 207 55 209 57
rect 203 54 209 55
rect 157 48 169 50
rect 157 46 162 48
rect 164 46 169 48
rect 157 44 169 46
rect 163 40 169 44
rect 163 38 164 40
rect 166 38 169 40
rect 163 36 169 38
rect 180 39 195 41
rect 180 37 186 39
rect 188 38 195 39
rect 188 37 191 38
rect 180 36 191 37
rect 193 36 195 38
rect 180 35 195 36
rect 180 29 186 35
rect 205 25 209 54
rect 68 16 77 17
rect 79 16 81 18
rect 68 13 81 16
rect 85 22 98 25
rect 85 20 87 22
rect 89 21 98 22
rect 132 23 145 25
rect 132 21 141 23
rect 143 21 145 23
rect 89 20 90 21
rect 139 20 145 21
rect 149 22 162 25
rect 149 20 151 22
rect 153 21 162 22
rect 196 23 209 25
rect 196 21 205 23
rect 207 21 209 23
rect 153 20 154 21
rect 203 20 209 21
rect 213 57 219 58
rect 213 55 215 57
rect 217 55 219 57
rect 213 54 219 55
rect 213 39 217 54
rect 213 37 214 39
rect 216 37 217 39
rect 213 25 217 37
rect 227 39 242 41
rect 227 38 234 39
rect 227 36 229 38
rect 231 37 234 38
rect 236 37 242 39
rect 231 36 242 37
rect 227 35 242 36
rect 236 29 242 35
rect 253 48 265 50
rect 253 46 257 48
rect 259 46 265 48
rect 253 44 265 46
rect 253 40 259 44
rect 253 38 256 40
rect 258 38 259 40
rect 253 36 259 38
rect 287 51 296 52
rect 287 49 289 51
rect 291 49 296 51
rect 287 48 296 49
rect 292 43 296 48
rect 276 42 288 43
rect 276 40 283 42
rect 285 40 288 42
rect 276 37 288 40
rect 292 39 304 43
rect 276 32 280 37
rect 300 36 304 39
rect 276 30 277 32
rect 279 30 280 32
rect 292 33 296 35
rect 292 31 293 33
rect 295 31 296 33
rect 292 30 296 31
rect 276 29 280 30
rect 284 26 296 30
rect 300 34 301 36
rect 303 34 304 36
rect 213 23 226 25
rect 213 21 215 23
rect 217 21 226 23
rect 260 22 273 25
rect 260 21 269 22
rect 213 20 219 21
rect 268 20 269 21
rect 271 20 273 22
rect 284 24 288 26
rect 284 22 285 24
rect 287 22 288 24
rect 284 21 288 22
rect 85 17 90 20
rect 149 18 154 20
rect 85 15 86 17
rect 88 15 90 17
rect 85 12 90 15
rect 81 7 85 8
rect 149 16 150 18
rect 152 16 154 18
rect 149 12 154 16
rect 268 17 273 20
rect 268 15 270 17
rect 272 15 273 17
rect 268 13 273 15
rect 300 17 304 34
rect 368 58 374 59
rect 368 56 370 58
rect 372 56 374 58
rect 368 55 374 56
rect 322 50 334 51
rect 322 48 326 50
rect 328 48 334 50
rect 322 45 334 48
rect 328 41 334 45
rect 328 39 329 41
rect 331 39 334 41
rect 328 37 334 39
rect 345 39 360 42
rect 345 37 347 39
rect 349 37 356 39
rect 358 37 360 39
rect 345 36 360 37
rect 345 30 351 36
rect 370 26 374 55
rect 422 57 444 58
rect 422 55 425 57
rect 427 55 444 57
rect 422 54 444 55
rect 502 57 507 59
rect 502 55 503 57
rect 505 55 507 57
rect 295 16 304 17
rect 295 14 297 16
rect 299 14 304 16
rect 295 13 304 14
rect 314 23 327 26
rect 314 21 316 23
rect 318 22 327 23
rect 361 24 374 26
rect 361 22 370 24
rect 372 22 374 24
rect 318 21 319 22
rect 368 21 374 22
rect 382 50 387 52
rect 382 48 384 50
rect 386 48 387 50
rect 382 46 387 48
rect 414 50 418 51
rect 414 48 415 50
rect 417 48 418 50
rect 382 39 386 46
rect 382 37 383 39
rect 385 37 386 39
rect 382 27 386 37
rect 414 42 418 48
rect 382 25 384 27
rect 314 17 319 21
rect 382 20 386 25
rect 314 15 316 17
rect 318 15 319 17
rect 314 13 319 15
rect 382 18 384 20
rect 397 41 418 42
rect 397 39 401 41
rect 403 39 418 41
rect 397 38 418 39
rect 422 34 426 54
rect 397 32 411 34
rect 413 32 418 34
rect 397 30 418 32
rect 414 28 418 30
rect 422 32 428 34
rect 422 30 425 32
rect 427 30 428 32
rect 422 28 428 30
rect 414 25 428 28
rect 414 24 425 25
rect 414 21 418 24
rect 422 23 425 24
rect 427 23 428 25
rect 422 21 428 23
rect 455 42 459 51
rect 502 53 507 55
rect 446 41 461 42
rect 446 39 450 41
rect 452 39 457 41
rect 459 39 461 41
rect 446 38 461 39
rect 471 41 479 43
rect 471 39 472 41
rect 474 39 476 41
rect 478 39 479 41
rect 471 37 479 39
rect 471 34 476 37
rect 438 30 476 34
rect 503 33 507 53
rect 503 31 504 33
rect 506 31 507 33
rect 502 29 507 31
rect 502 27 503 29
rect 505 27 507 29
rect 502 22 507 27
rect 502 20 503 22
rect 505 20 507 22
rect 511 57 533 58
rect 511 55 514 57
rect 516 55 533 57
rect 511 54 533 55
rect 591 57 596 59
rect 591 55 592 57
rect 594 55 596 57
rect 511 50 515 54
rect 511 48 512 50
rect 514 48 515 50
rect 511 34 515 48
rect 544 50 548 51
rect 544 48 545 50
rect 547 48 548 50
rect 511 32 517 34
rect 511 30 514 32
rect 516 30 517 32
rect 511 25 517 30
rect 511 23 514 25
rect 516 23 517 25
rect 511 21 517 23
rect 544 42 548 48
rect 591 53 596 55
rect 592 51 593 53
rect 595 51 596 53
rect 535 41 550 42
rect 535 39 539 41
rect 541 39 546 41
rect 548 39 550 41
rect 535 38 550 39
rect 560 41 568 43
rect 560 39 565 41
rect 567 39 568 41
rect 560 37 568 39
rect 560 34 565 37
rect 527 33 565 34
rect 527 31 534 33
rect 536 31 565 33
rect 527 30 565 31
rect 592 31 596 51
rect 591 29 596 31
rect 656 57 660 59
rect 655 55 660 57
rect 655 53 656 55
rect 658 53 660 55
rect 655 51 660 53
rect 607 49 620 50
rect 607 47 617 49
rect 619 47 620 49
rect 607 46 620 47
rect 614 41 620 46
rect 614 39 615 41
rect 617 39 620 41
rect 614 37 620 39
rect 640 36 644 43
rect 640 35 642 36
rect 632 34 642 35
rect 632 33 644 34
rect 632 31 637 33
rect 639 31 644 33
rect 632 29 644 31
rect 591 27 592 29
rect 594 27 596 29
rect 591 22 596 27
rect 502 18 507 20
rect 591 20 592 22
rect 594 20 596 22
rect 591 18 596 20
rect 382 14 395 18
rect 382 13 386 14
rect 494 14 507 18
rect 583 14 596 18
rect 600 22 613 26
rect 600 21 605 22
rect 656 41 660 51
rect 656 39 657 41
rect 659 39 660 41
rect 600 19 602 21
rect 604 19 605 21
rect 600 18 605 19
rect 600 16 602 18
rect 604 16 605 18
rect 656 18 660 39
rect 664 50 668 59
rect 664 48 666 50
rect 664 46 668 48
rect 664 44 665 46
rect 667 44 668 46
rect 664 32 668 44
rect 672 43 676 51
rect 672 41 684 43
rect 672 39 673 41
rect 675 39 680 41
rect 682 39 684 41
rect 672 37 684 39
rect 664 30 666 32
rect 664 27 668 30
rect 664 25 676 27
rect 664 23 666 25
rect 668 23 676 25
rect 664 21 676 23
rect 647 17 660 18
rect 600 13 605 16
rect 647 15 656 17
rect 658 15 660 17
rect 647 14 660 15
rect 276 7 688 8
rect -18 6 317 7
rect -18 4 7 6
rect 9 4 21 6
rect 23 4 35 6
rect 37 4 76 6
rect 78 4 88 6
rect 90 4 152 6
rect 154 4 268 6
rect 270 5 317 6
rect 319 5 385 7
rect 387 5 667 7
rect 669 5 679 7
rect 681 5 688 7
rect 270 4 688 5
rect -18 0 688 4
rect -18 -1 -11 0
<< alu2 >>
rect 524 282 547 286
rect 369 278 374 280
rect 524 279 528 282
rect 369 276 370 278
rect 372 276 374 278
rect 4 262 52 263
rect 4 260 49 262
rect 51 260 52 262
rect 4 259 52 260
rect 151 262 185 263
rect 151 260 152 262
rect 154 260 182 262
rect 184 260 185 262
rect 151 259 185 260
rect 4 254 9 259
rect 302 256 343 257
rect 4 252 6 254
rect 8 252 9 254
rect 4 189 9 252
rect 28 254 217 255
rect 28 252 29 254
rect 31 252 214 254
rect 216 252 217 254
rect 302 254 303 256
rect 305 254 339 256
rect 341 254 343 256
rect 302 253 343 254
rect 28 251 217 252
rect 20 249 24 250
rect 20 247 21 249
rect 23 247 24 249
rect 20 246 72 247
rect 20 244 69 246
rect 71 244 72 246
rect 20 243 72 244
rect 140 245 144 247
rect 140 243 141 245
rect 143 243 144 245
rect 92 242 96 243
rect 92 240 93 242
rect 95 240 96 242
rect 92 229 96 240
rect 140 238 144 243
rect 173 245 364 246
rect 173 243 174 245
rect 176 243 178 245
rect 180 243 271 245
rect 273 243 360 245
rect 362 243 364 245
rect 173 242 364 243
rect 140 234 265 238
rect 92 225 232 229
rect 36 196 97 197
rect 36 194 37 196
rect 39 194 94 196
rect 96 194 97 196
rect 36 193 97 194
rect 141 195 169 197
rect 141 193 142 195
rect 144 193 162 195
rect 164 193 169 195
rect 141 191 169 193
rect 4 187 49 189
rect 227 188 232 225
rect 259 197 265 234
rect 369 228 374 276
rect 400 278 528 279
rect 543 279 547 282
rect 543 278 603 279
rect 400 276 416 278
rect 418 276 472 278
rect 474 276 528 278
rect 400 275 528 276
rect 533 277 539 278
rect 533 275 536 277
rect 538 275 539 277
rect 543 276 600 278
rect 602 276 603 278
rect 543 275 603 276
rect 400 271 404 275
rect 533 271 539 275
rect 400 269 401 271
rect 403 269 404 271
rect 400 268 404 269
rect 408 270 539 271
rect 408 268 535 270
rect 537 268 539 270
rect 408 267 539 268
rect 630 272 669 273
rect 630 270 632 272
rect 634 270 665 272
rect 667 270 669 272
rect 630 269 669 270
rect 408 263 412 267
rect 630 264 635 269
rect 300 223 374 228
rect 384 259 388 262
rect 408 261 409 263
rect 411 261 412 263
rect 408 259 412 261
rect 622 263 635 264
rect 622 261 623 263
rect 625 261 635 263
rect 622 260 635 261
rect 567 259 611 260
rect 384 257 385 259
rect 387 257 388 259
rect 253 195 271 197
rect 253 193 257 195
rect 259 193 271 195
rect 253 191 271 193
rect 4 185 5 187
rect 7 185 46 187
rect 48 185 49 187
rect 4 183 49 185
rect 180 186 217 188
rect 180 184 186 186
rect 188 184 214 186
rect 216 184 217 186
rect 77 183 121 184
rect 77 181 78 183
rect 80 181 117 183
rect 119 181 121 183
rect 180 182 217 184
rect 227 186 239 188
rect 227 184 234 186
rect 236 184 239 186
rect 227 182 239 184
rect 300 183 304 223
rect 384 218 388 257
rect 449 256 461 258
rect 449 254 452 256
rect 454 254 461 256
rect 449 252 461 254
rect 471 256 508 258
rect 567 257 569 259
rect 571 257 608 259
rect 610 257 611 259
rect 567 256 611 257
rect 471 254 472 256
rect 474 254 500 256
rect 502 254 508 256
rect 471 252 508 254
rect 639 255 684 257
rect 639 253 640 255
rect 642 253 681 255
rect 683 253 684 255
rect 417 247 435 249
rect 417 245 429 247
rect 431 245 435 247
rect 417 243 435 245
rect 300 181 301 183
rect 303 181 304 183
rect 77 180 121 181
rect 53 179 66 180
rect 53 177 63 179
rect 65 177 66 179
rect 53 176 66 177
rect 276 179 280 181
rect 276 177 277 179
rect 279 177 280 179
rect 300 178 304 181
rect 314 213 388 218
rect 53 171 58 176
rect 276 173 280 177
rect 19 170 58 171
rect 19 168 21 170
rect 23 168 54 170
rect 56 168 58 170
rect 19 167 58 168
rect 149 169 280 173
rect 284 171 288 172
rect 284 169 285 171
rect 287 169 288 171
rect 149 165 155 169
rect 284 165 288 169
rect 85 164 145 165
rect 85 162 86 164
rect 88 162 145 164
rect 149 163 150 165
rect 152 163 155 165
rect 149 162 155 163
rect 160 164 288 165
rect 160 162 270 164
rect 272 162 288 164
rect 85 161 145 162
rect 141 158 145 161
rect 160 161 288 162
rect 314 164 319 213
rect 423 206 429 243
rect 456 215 461 252
rect 639 251 684 253
rect 519 247 547 249
rect 519 245 524 247
rect 526 245 544 247
rect 546 245 547 247
rect 519 243 547 245
rect 591 246 652 247
rect 591 244 592 246
rect 594 244 649 246
rect 651 244 652 246
rect 591 243 652 244
rect 456 211 596 215
rect 423 204 548 206
rect 423 202 545 204
rect 547 202 548 204
rect 324 197 515 198
rect 324 195 326 197
rect 328 195 415 197
rect 417 195 508 197
rect 510 195 512 197
rect 514 195 515 197
rect 324 194 515 195
rect 544 197 548 202
rect 592 200 596 211
rect 592 198 593 200
rect 595 198 596 200
rect 592 197 596 198
rect 544 195 545 197
rect 547 195 548 197
rect 544 193 548 195
rect 616 196 668 197
rect 616 194 617 196
rect 619 194 668 196
rect 616 193 668 194
rect 664 191 665 193
rect 667 191 668 193
rect 664 190 668 191
rect 471 188 660 189
rect 345 186 386 187
rect 345 184 347 186
rect 349 184 383 186
rect 385 184 386 186
rect 471 186 472 188
rect 474 186 657 188
rect 659 186 660 188
rect 471 185 660 186
rect 679 188 684 251
rect 679 186 680 188
rect 682 186 684 188
rect 345 183 386 184
rect 679 181 684 186
rect 503 180 537 181
rect 370 178 381 179
rect 370 176 371 178
rect 373 176 377 178
rect 379 176 381 178
rect 503 178 504 180
rect 506 178 534 180
rect 536 178 537 180
rect 503 177 537 178
rect 636 180 684 181
rect 636 178 637 180
rect 639 178 684 180
rect 636 177 684 178
rect 370 174 381 176
rect 600 171 605 173
rect 600 169 602 171
rect 604 169 605 171
rect 600 164 605 169
rect 314 162 316 164
rect 318 162 319 164
rect 160 158 164 161
rect 314 160 319 162
rect 597 163 605 164
rect 597 161 602 163
rect 604 161 605 163
rect 597 160 605 161
rect 141 154 164 158
rect 524 135 547 139
rect 369 131 374 133
rect 524 132 528 135
rect 369 129 370 131
rect 372 129 374 131
rect 4 115 52 116
rect 4 113 49 115
rect 51 113 52 115
rect 4 112 52 113
rect 151 115 185 116
rect 151 113 152 115
rect 154 113 182 115
rect 184 113 185 115
rect 151 112 185 113
rect 4 107 9 112
rect 302 109 343 110
rect 4 105 6 107
rect 8 105 9 107
rect 4 42 9 105
rect 28 107 217 108
rect 28 105 29 107
rect 31 105 214 107
rect 216 105 217 107
rect 302 107 303 109
rect 305 107 339 109
rect 341 107 343 109
rect 302 106 343 107
rect 28 104 217 105
rect 20 102 24 103
rect 20 100 21 102
rect 23 100 24 102
rect 20 99 72 100
rect 20 97 69 99
rect 71 97 72 99
rect 20 96 72 97
rect 140 98 144 100
rect 140 96 141 98
rect 143 96 144 98
rect 92 95 96 96
rect 92 93 93 95
rect 95 93 96 95
rect 92 82 96 93
rect 140 91 144 96
rect 173 98 364 99
rect 173 96 174 98
rect 176 96 178 98
rect 180 96 271 98
rect 273 96 360 98
rect 362 96 364 98
rect 173 95 364 96
rect 140 87 265 91
rect 92 78 232 82
rect 36 49 97 50
rect 36 47 37 49
rect 39 47 94 49
rect 96 47 97 49
rect 36 46 97 47
rect 141 48 169 50
rect 141 46 142 48
rect 144 46 162 48
rect 164 46 169 48
rect 141 44 169 46
rect 4 40 49 42
rect 227 41 232 78
rect 259 50 265 87
rect 369 80 374 129
rect 400 131 528 132
rect 543 132 547 135
rect 543 131 603 132
rect 400 129 416 131
rect 418 129 471 131
rect 473 129 528 131
rect 400 128 528 129
rect 533 130 539 131
rect 533 128 536 130
rect 538 128 539 130
rect 543 129 600 131
rect 602 129 603 131
rect 543 128 603 129
rect 400 124 404 128
rect 533 124 539 128
rect 400 122 401 124
rect 403 122 404 124
rect 400 121 404 122
rect 408 123 539 124
rect 408 121 535 123
rect 537 121 539 123
rect 408 120 539 121
rect 630 125 669 126
rect 630 123 632 125
rect 634 123 665 125
rect 667 123 669 125
rect 630 122 669 123
rect 408 116 412 120
rect 630 117 635 122
rect 300 75 374 80
rect 384 112 388 115
rect 408 114 409 116
rect 411 114 412 116
rect 408 112 412 114
rect 622 116 635 117
rect 622 114 623 116
rect 625 114 635 116
rect 622 113 635 114
rect 567 112 611 113
rect 384 110 385 112
rect 387 110 388 112
rect 253 48 271 50
rect 253 46 257 48
rect 259 46 271 48
rect 253 44 271 46
rect 4 38 5 40
rect 7 38 46 40
rect 48 38 49 40
rect 4 36 49 38
rect 180 39 217 41
rect 180 37 186 39
rect 188 37 214 39
rect 216 37 217 39
rect 77 36 121 37
rect 77 34 78 36
rect 80 34 117 36
rect 119 34 121 36
rect 180 35 217 37
rect 227 39 239 41
rect 227 37 234 39
rect 236 37 239 39
rect 227 35 239 37
rect 300 36 304 75
rect 384 70 388 110
rect 449 109 461 111
rect 449 107 452 109
rect 454 107 461 109
rect 449 105 461 107
rect 471 109 508 111
rect 567 110 569 112
rect 571 110 608 112
rect 610 110 611 112
rect 567 109 611 110
rect 471 107 472 109
rect 474 107 500 109
rect 502 107 508 109
rect 471 105 508 107
rect 639 108 684 110
rect 639 106 640 108
rect 642 106 681 108
rect 683 106 684 108
rect 417 100 435 102
rect 417 98 424 100
rect 426 98 429 100
rect 431 98 435 100
rect 417 96 435 98
rect 300 34 301 36
rect 303 34 304 36
rect 77 33 121 34
rect 53 32 66 33
rect 53 30 63 32
rect 65 30 66 32
rect 53 29 66 30
rect 276 32 280 34
rect 276 30 277 32
rect 279 30 280 32
rect 300 31 304 34
rect 314 65 388 70
rect 53 24 58 29
rect 276 26 280 30
rect 19 23 58 24
rect 19 21 21 23
rect 23 21 54 23
rect 56 21 58 23
rect 19 20 58 21
rect 149 22 280 26
rect 284 24 288 25
rect 284 22 285 24
rect 287 22 288 24
rect 149 18 155 22
rect 284 18 288 22
rect 85 17 145 18
rect 85 15 86 17
rect 88 15 145 17
rect 149 16 150 18
rect 152 16 155 18
rect 149 15 155 16
rect 160 17 288 18
rect 160 15 270 17
rect 272 15 288 17
rect 85 14 145 15
rect 141 11 145 14
rect 160 14 288 15
rect 314 17 319 65
rect 423 59 429 96
rect 456 68 461 105
rect 639 104 684 106
rect 519 100 547 102
rect 519 98 524 100
rect 526 98 544 100
rect 546 98 547 100
rect 519 96 547 98
rect 591 99 652 100
rect 591 97 592 99
rect 594 97 649 99
rect 651 97 652 99
rect 591 96 652 97
rect 456 64 596 68
rect 423 55 548 59
rect 324 50 515 51
rect 324 48 326 50
rect 328 48 415 50
rect 417 48 508 50
rect 510 48 512 50
rect 514 48 515 50
rect 324 47 515 48
rect 544 50 548 55
rect 592 53 596 64
rect 592 51 593 53
rect 595 51 596 53
rect 592 50 596 51
rect 544 48 545 50
rect 547 48 548 50
rect 544 46 548 48
rect 616 49 668 50
rect 616 47 617 49
rect 619 47 668 49
rect 616 46 668 47
rect 664 44 665 46
rect 667 44 668 46
rect 664 43 668 44
rect 471 41 660 42
rect 345 39 386 40
rect 345 37 347 39
rect 349 37 383 39
rect 385 37 386 39
rect 471 39 472 41
rect 474 39 657 41
rect 659 39 660 41
rect 471 38 660 39
rect 679 41 684 104
rect 679 39 680 41
rect 682 39 684 41
rect 345 36 386 37
rect 679 34 684 39
rect 503 33 537 34
rect 503 31 504 33
rect 506 31 534 33
rect 536 31 537 33
rect 503 30 537 31
rect 636 33 684 34
rect 636 31 637 33
rect 639 31 684 33
rect 636 30 684 31
rect 314 15 316 17
rect 318 15 319 17
rect 160 11 164 14
rect 314 13 319 15
rect 600 24 612 26
rect 600 22 602 24
rect 604 22 612 24
rect 600 18 605 22
rect 600 16 602 18
rect 604 16 605 18
rect 600 15 605 16
rect 600 13 602 15
rect 604 13 605 15
rect 600 12 605 13
rect 141 7 164 11
<< alu3 >>
rect 534 280 539 281
rect 471 278 481 279
rect 471 276 472 278
rect 474 276 476 278
rect 478 276 481 278
rect 471 275 481 276
rect 534 278 536 280
rect 538 278 539 280
rect 534 270 539 278
rect 534 268 535 270
rect 537 268 539 270
rect 534 267 539 268
rect 622 263 626 264
rect 622 261 623 263
rect 625 261 626 263
rect 177 245 181 246
rect 177 243 178 245
rect 180 243 181 245
rect 177 222 181 243
rect 622 222 626 261
rect 62 218 181 222
rect 507 218 626 222
rect 62 179 66 218
rect 507 197 511 218
rect 507 195 508 197
rect 510 195 511 197
rect 507 194 511 195
rect 544 204 548 206
rect 544 202 545 204
rect 547 202 548 204
rect 62 177 63 179
rect 65 177 66 179
rect 62 176 66 177
rect 376 178 381 179
rect 376 176 377 178
rect 379 176 381 178
rect 376 160 381 176
rect 544 164 548 202
rect 600 164 605 173
rect 544 163 605 164
rect 544 161 598 163
rect 600 161 602 163
rect 604 161 605 163
rect 544 160 605 161
rect 376 155 428 160
rect 423 100 428 155
rect 534 133 539 135
rect 468 131 479 132
rect 468 129 471 131
rect 473 129 476 131
rect 478 129 479 131
rect 468 128 479 129
rect 534 131 536 133
rect 538 131 539 133
rect 534 124 539 131
rect 526 123 539 124
rect 526 121 535 123
rect 537 121 539 123
rect 526 120 539 121
rect 177 98 181 99
rect 177 96 178 98
rect 180 96 181 98
rect 423 98 424 100
rect 426 98 428 100
rect 423 96 428 98
rect 622 116 626 117
rect 622 114 623 116
rect 625 114 626 116
rect 177 75 181 96
rect 622 75 626 114
rect 62 71 181 75
rect 507 71 626 75
rect 62 32 66 71
rect 507 50 511 71
rect 507 48 508 50
rect 510 48 511 50
rect 507 47 511 48
rect 62 30 63 32
rect 65 30 66 32
rect 62 29 66 30
rect 600 25 612 26
rect 600 24 606 25
rect 600 22 602 24
rect 604 23 606 24
rect 608 23 612 25
rect 604 22 612 23
rect 600 15 605 22
rect 600 13 602 15
rect 604 13 605 15
rect 600 12 605 13
<< alu4 >>
rect 534 280 539 281
rect 475 278 479 279
rect 475 276 476 278
rect 478 276 479 278
rect 36 192 40 196
rect 475 131 479 276
rect 475 129 476 131
rect 478 129 479 131
rect 475 128 479 129
rect 534 278 536 280
rect 538 278 539 280
rect 534 133 539 278
rect 648 244 652 248
rect 600 164 605 173
rect 596 163 605 164
rect 596 161 598 163
rect 600 161 605 163
rect 596 160 605 161
rect 534 131 536 133
rect 538 131 539 133
rect 534 120 539 131
rect 36 45 40 49
rect 600 26 605 160
rect 648 97 652 101
rect 600 25 612 26
rect 600 23 606 25
rect 608 23 612 25
rect 600 22 612 23
rect 600 12 605 22
<< ptie >>
rect 5 228 23 230
rect 5 226 7 228
rect 9 226 19 228
rect 21 226 23 228
rect 5 224 23 226
rect 299 228 305 230
rect 299 226 301 228
rect 303 226 305 228
rect 299 224 305 226
rect 385 228 411 230
rect 385 226 387 228
rect 389 226 407 228
rect 409 226 411 228
rect 385 224 411 226
rect 608 229 642 231
rect 608 227 610 229
rect 612 227 638 229
rect 640 227 642 229
rect 608 225 642 227
rect 649 229 655 231
rect 649 227 651 229
rect 653 227 655 229
rect 649 225 655 227
rect 33 213 39 215
rect 33 211 35 213
rect 37 211 39 213
rect 33 209 39 211
rect 46 213 80 215
rect 46 211 48 213
rect 50 211 76 213
rect 78 211 80 213
rect 46 209 80 211
rect 277 214 303 216
rect 277 212 279 214
rect 281 212 299 214
rect 301 212 303 214
rect 277 210 303 212
rect 383 214 389 216
rect 383 212 385 214
rect 387 212 389 214
rect 383 210 389 212
rect 665 214 683 216
rect 665 212 667 214
rect 669 212 679 214
rect 681 212 683 214
rect 665 210 683 212
rect 5 81 23 83
rect 5 79 7 81
rect 9 79 19 81
rect 21 79 23 81
rect 5 77 23 79
rect 299 81 305 83
rect 299 79 301 81
rect 303 79 305 81
rect 299 77 305 79
rect 385 81 411 83
rect 385 79 387 81
rect 389 79 407 81
rect 409 79 411 81
rect 385 77 411 79
rect 608 82 642 84
rect 608 80 610 82
rect 612 80 638 82
rect 640 80 642 82
rect 608 78 642 80
rect 649 82 655 84
rect 649 80 651 82
rect 653 80 655 82
rect 649 78 655 80
rect 33 66 39 68
rect 33 64 35 66
rect 37 64 39 66
rect 33 62 39 64
rect 46 66 80 68
rect 46 64 48 66
rect 50 64 76 66
rect 78 64 80 66
rect 46 62 80 64
rect 277 67 303 69
rect 277 65 279 67
rect 281 65 299 67
rect 301 65 303 67
rect 277 63 303 65
rect 383 67 389 69
rect 383 65 385 67
rect 387 65 389 67
rect 383 63 389 65
rect 665 67 683 69
rect 665 65 667 67
rect 669 65 679 67
rect 681 65 683 67
rect 665 63 683 65
<< ntie >>
rect 5 288 23 290
rect 5 286 7 288
rect 9 286 19 288
rect 21 286 23 288
rect 5 284 23 286
rect 299 288 305 290
rect 299 286 301 288
rect 303 286 305 288
rect 299 284 305 286
rect 367 288 373 290
rect 367 286 369 288
rect 371 286 373 288
rect 416 289 422 291
rect 416 287 418 289
rect 420 287 422 289
rect 367 284 373 286
rect 416 285 422 287
rect 532 289 538 291
rect 532 287 534 289
rect 536 287 538 289
rect 532 285 538 287
rect 596 289 602 291
rect 596 287 598 289
rect 600 287 602 289
rect 596 285 602 287
rect 608 289 614 291
rect 608 287 610 289
rect 612 287 614 289
rect 649 289 683 291
rect 608 285 614 287
rect 649 287 651 289
rect 653 287 665 289
rect 667 287 679 289
rect 681 287 683 289
rect 649 285 683 287
rect 5 153 39 155
rect 5 151 7 153
rect 9 151 21 153
rect 23 151 35 153
rect 37 151 39 153
rect 74 153 80 155
rect 5 149 39 151
rect 74 151 76 153
rect 78 151 80 153
rect 74 149 80 151
rect 86 153 92 155
rect 86 151 88 153
rect 90 151 92 153
rect 86 149 92 151
rect 150 153 156 155
rect 150 151 152 153
rect 154 151 156 153
rect 150 149 156 151
rect 266 153 272 155
rect 315 154 321 156
rect 266 151 268 153
rect 270 151 272 153
rect 266 149 272 151
rect 315 152 317 154
rect 319 152 321 154
rect 315 150 321 152
rect 383 154 389 156
rect 383 152 385 154
rect 387 152 389 154
rect 383 150 389 152
rect 665 154 683 156
rect 665 152 667 154
rect 669 152 679 154
rect 681 152 683 154
rect 665 150 683 152
rect 5 141 23 143
rect 5 139 7 141
rect 9 139 19 141
rect 21 139 23 141
rect 5 137 23 139
rect 299 141 305 143
rect 299 139 301 141
rect 303 139 305 141
rect 299 137 305 139
rect 367 141 373 143
rect 367 139 369 141
rect 371 139 373 141
rect 416 142 422 144
rect 416 140 418 142
rect 420 140 422 142
rect 367 137 373 139
rect 416 138 422 140
rect 532 142 538 144
rect 532 140 534 142
rect 536 140 538 142
rect 532 138 538 140
rect 596 142 602 144
rect 596 140 598 142
rect 600 140 602 142
rect 596 138 602 140
rect 608 142 614 144
rect 608 140 610 142
rect 612 140 614 142
rect 649 142 683 144
rect 608 138 614 140
rect 649 140 651 142
rect 653 140 665 142
rect 667 140 679 142
rect 681 140 683 142
rect 649 138 683 140
rect 5 6 39 8
rect 5 4 7 6
rect 9 4 21 6
rect 23 4 35 6
rect 37 4 39 6
rect 74 6 80 8
rect 5 2 39 4
rect 74 4 76 6
rect 78 4 80 6
rect 74 2 80 4
rect 86 6 92 8
rect 86 4 88 6
rect 90 4 92 6
rect 86 2 92 4
rect 150 6 156 8
rect 150 4 152 6
rect 154 4 156 6
rect 150 2 156 4
rect 266 6 272 8
rect 315 7 321 9
rect 266 4 268 6
rect 270 4 272 6
rect 266 2 272 4
rect 315 5 317 7
rect 319 5 321 7
rect 315 3 321 5
rect 383 7 389 9
rect 383 5 385 7
rect 387 5 389 7
rect 383 3 389 5
rect 665 7 683 9
rect 665 5 667 7
rect 669 5 679 7
rect 681 5 683 7
rect 665 3 683 5
<< nmos >>
rect 15 238 17 247
rect 35 233 37 242
rect 45 233 47 241
rect 52 233 54 241
rect 62 233 64 241
rect 69 233 71 241
rect 79 235 81 241
rect 99 227 101 240
rect 109 230 111 240
rect 119 233 121 247
rect 129 233 131 247
rect 149 227 151 247
rect 156 227 158 247
rect 167 227 169 241
rect 188 227 190 240
rect 198 230 200 240
rect 208 233 210 247
rect 218 233 220 247
rect 238 227 240 247
rect 245 227 247 247
rect 277 241 279 247
rect 287 241 289 247
rect 256 227 258 241
rect 297 238 299 247
rect 392 240 394 246
rect 402 240 404 246
rect 321 233 323 239
rect 331 233 333 239
rect 338 233 340 239
rect 348 233 350 239
rect 355 233 357 239
rect 365 233 367 239
rect 422 234 424 240
rect 432 234 434 240
rect 439 234 441 240
rect 449 234 451 240
rect 456 234 458 240
rect 466 234 468 240
rect 486 234 488 240
rect 496 234 498 240
rect 503 234 505 240
rect 513 234 515 240
rect 520 234 522 240
rect 530 234 532 240
rect 550 234 552 240
rect 560 234 562 240
rect 567 234 569 240
rect 577 234 579 240
rect 584 234 586 240
rect 594 234 596 240
rect 614 237 616 243
rect 624 237 626 243
rect 634 237 636 243
rect 655 237 657 243
rect 667 231 669 240
rect 674 231 676 240
rect 12 200 14 209
rect 19 200 21 209
rect 31 197 33 203
rect 52 197 54 203
rect 62 197 64 203
rect 72 197 74 203
rect 92 200 94 206
rect 102 200 104 206
rect 109 200 111 206
rect 119 200 121 206
rect 126 200 128 206
rect 136 200 138 206
rect 156 200 158 206
rect 166 200 168 206
rect 173 200 175 206
rect 183 200 185 206
rect 190 200 192 206
rect 200 200 202 206
rect 220 200 222 206
rect 230 200 232 206
rect 237 200 239 206
rect 247 200 249 206
rect 254 200 256 206
rect 264 200 266 206
rect 321 201 323 207
rect 331 201 333 207
rect 338 201 340 207
rect 348 201 350 207
rect 355 201 357 207
rect 365 201 367 207
rect 284 194 286 200
rect 294 194 296 200
rect 389 193 391 202
rect 430 199 432 213
rect 399 193 401 199
rect 409 193 411 199
rect 441 193 443 213
rect 448 193 450 213
rect 468 193 470 207
rect 478 193 480 207
rect 488 200 490 210
rect 498 200 500 213
rect 519 199 521 213
rect 530 193 532 213
rect 537 193 539 213
rect 557 193 559 207
rect 567 193 569 207
rect 577 200 579 210
rect 587 200 589 213
rect 607 199 609 205
rect 617 199 619 207
rect 624 199 626 207
rect 634 199 636 207
rect 641 199 643 207
rect 651 198 653 207
rect 671 193 673 202
rect 15 91 17 100
rect 35 86 37 95
rect 45 86 47 94
rect 52 86 54 94
rect 62 86 64 94
rect 69 86 71 94
rect 79 88 81 94
rect 99 80 101 93
rect 109 83 111 93
rect 119 86 121 100
rect 129 86 131 100
rect 149 80 151 100
rect 156 80 158 100
rect 167 80 169 94
rect 188 80 190 93
rect 198 83 200 93
rect 208 86 210 100
rect 218 86 220 100
rect 238 80 240 100
rect 245 80 247 100
rect 277 94 279 100
rect 287 94 289 100
rect 256 80 258 94
rect 297 91 299 100
rect 392 93 394 99
rect 402 93 404 99
rect 321 86 323 92
rect 331 86 333 92
rect 338 86 340 92
rect 348 86 350 92
rect 355 86 357 92
rect 365 86 367 92
rect 422 87 424 93
rect 432 87 434 93
rect 439 87 441 93
rect 449 87 451 93
rect 456 87 458 93
rect 466 87 468 93
rect 486 87 488 93
rect 496 87 498 93
rect 503 87 505 93
rect 513 87 515 93
rect 520 87 522 93
rect 530 87 532 93
rect 550 87 552 93
rect 560 87 562 93
rect 567 87 569 93
rect 577 87 579 93
rect 584 87 586 93
rect 594 87 596 93
rect 614 90 616 96
rect 624 90 626 96
rect 634 90 636 96
rect 655 90 657 96
rect 667 84 669 93
rect 674 84 676 93
rect 12 53 14 62
rect 19 53 21 62
rect 31 50 33 56
rect 52 50 54 56
rect 62 50 64 56
rect 72 50 74 56
rect 92 53 94 59
rect 102 53 104 59
rect 109 53 111 59
rect 119 53 121 59
rect 126 53 128 59
rect 136 53 138 59
rect 156 53 158 59
rect 166 53 168 59
rect 173 53 175 59
rect 183 53 185 59
rect 190 53 192 59
rect 200 53 202 59
rect 220 53 222 59
rect 230 53 232 59
rect 237 53 239 59
rect 247 53 249 59
rect 254 53 256 59
rect 264 53 266 59
rect 321 54 323 60
rect 331 54 333 60
rect 338 54 340 60
rect 348 54 350 60
rect 355 54 357 60
rect 365 54 367 60
rect 284 47 286 53
rect 294 47 296 53
rect 389 46 391 55
rect 430 52 432 66
rect 399 46 401 52
rect 409 46 411 52
rect 441 46 443 66
rect 448 46 450 66
rect 468 46 470 60
rect 478 46 480 60
rect 488 53 490 63
rect 498 53 500 66
rect 519 52 521 66
rect 530 46 532 66
rect 537 46 539 66
rect 557 46 559 60
rect 567 46 569 60
rect 577 53 579 63
rect 587 53 589 66
rect 607 52 609 58
rect 617 52 619 60
rect 624 52 626 60
rect 634 52 636 60
rect 641 52 643 60
rect 651 51 653 60
rect 671 46 673 55
<< pmos >>
rect 15 259 17 277
rect 35 269 37 287
rect 45 271 47 287
rect 52 271 54 287
rect 62 271 64 287
rect 69 271 71 287
rect 79 259 81 267
rect 99 262 101 287
rect 112 262 114 275
rect 122 259 124 284
rect 129 259 131 284
rect 147 259 149 287
rect 157 259 159 287
rect 167 259 169 287
rect 188 262 190 287
rect 201 262 203 275
rect 211 259 213 284
rect 218 259 220 284
rect 236 259 238 287
rect 246 259 248 287
rect 256 259 258 287
rect 277 266 279 287
rect 284 266 286 287
rect 297 259 299 277
rect 321 267 323 279
rect 331 267 333 279
rect 338 267 340 279
rect 348 267 350 279
rect 355 267 357 279
rect 394 267 396 287
rect 401 267 403 287
rect 365 259 367 265
rect 432 268 434 280
rect 439 268 441 280
rect 449 268 451 280
rect 456 268 458 280
rect 466 268 468 280
rect 486 268 488 280
rect 496 268 498 280
rect 503 268 505 280
rect 513 268 515 280
rect 520 268 522 280
rect 422 260 424 266
rect 550 268 552 280
rect 560 268 562 280
rect 567 268 569 280
rect 577 268 579 280
rect 584 268 586 280
rect 530 260 532 266
rect 614 267 616 279
rect 627 270 629 288
rect 634 270 636 288
rect 594 260 596 266
rect 655 260 657 272
rect 665 260 667 270
rect 675 260 677 270
rect 11 170 13 180
rect 21 170 23 180
rect 31 168 33 180
rect 92 174 94 180
rect 52 152 54 170
rect 59 152 61 170
rect 72 161 74 173
rect 156 174 158 180
rect 102 160 104 172
rect 109 160 111 172
rect 119 160 121 172
rect 126 160 128 172
rect 136 160 138 172
rect 264 174 266 180
rect 166 160 168 172
rect 173 160 175 172
rect 183 160 185 172
rect 190 160 192 172
rect 200 160 202 172
rect 220 160 222 172
rect 230 160 232 172
rect 237 160 239 172
rect 247 160 249 172
rect 254 160 256 172
rect 321 175 323 181
rect 285 153 287 173
rect 292 153 294 173
rect 331 161 333 173
rect 338 161 340 173
rect 348 161 350 173
rect 355 161 357 173
rect 365 161 367 173
rect 389 163 391 181
rect 402 153 404 174
rect 409 153 411 174
rect 430 153 432 181
rect 440 153 442 181
rect 450 153 452 181
rect 468 156 470 181
rect 475 156 477 181
rect 485 165 487 178
rect 498 153 500 178
rect 519 153 521 181
rect 529 153 531 181
rect 539 153 541 181
rect 557 156 559 181
rect 564 156 566 181
rect 574 165 576 178
rect 587 153 589 178
rect 607 173 609 181
rect 617 153 619 169
rect 624 153 626 169
rect 634 153 636 169
rect 641 153 643 169
rect 651 153 653 171
rect 671 163 673 181
rect 15 112 17 130
rect 35 122 37 140
rect 45 124 47 140
rect 52 124 54 140
rect 62 124 64 140
rect 69 124 71 140
rect 79 112 81 120
rect 99 115 101 140
rect 112 115 114 128
rect 122 112 124 137
rect 129 112 131 137
rect 147 112 149 140
rect 157 112 159 140
rect 167 112 169 140
rect 188 115 190 140
rect 201 115 203 128
rect 211 112 213 137
rect 218 112 220 137
rect 236 112 238 140
rect 246 112 248 140
rect 256 112 258 140
rect 277 119 279 140
rect 284 119 286 140
rect 297 112 299 130
rect 321 120 323 132
rect 331 120 333 132
rect 338 120 340 132
rect 348 120 350 132
rect 355 120 357 132
rect 394 120 396 140
rect 401 120 403 140
rect 365 112 367 118
rect 432 121 434 133
rect 439 121 441 133
rect 449 121 451 133
rect 456 121 458 133
rect 466 121 468 133
rect 486 121 488 133
rect 496 121 498 133
rect 503 121 505 133
rect 513 121 515 133
rect 520 121 522 133
rect 422 113 424 119
rect 550 121 552 133
rect 560 121 562 133
rect 567 121 569 133
rect 577 121 579 133
rect 584 121 586 133
rect 530 113 532 119
rect 614 120 616 132
rect 627 123 629 141
rect 634 123 636 141
rect 594 113 596 119
rect 655 113 657 125
rect 665 113 667 123
rect 675 113 677 123
rect 11 23 13 33
rect 21 23 23 33
rect 31 21 33 33
rect 92 27 94 33
rect 52 5 54 23
rect 59 5 61 23
rect 72 14 74 26
rect 156 27 158 33
rect 102 13 104 25
rect 109 13 111 25
rect 119 13 121 25
rect 126 13 128 25
rect 136 13 138 25
rect 264 27 266 33
rect 166 13 168 25
rect 173 13 175 25
rect 183 13 185 25
rect 190 13 192 25
rect 200 13 202 25
rect 220 13 222 25
rect 230 13 232 25
rect 237 13 239 25
rect 247 13 249 25
rect 254 13 256 25
rect 321 28 323 34
rect 285 6 287 26
rect 292 6 294 26
rect 331 14 333 26
rect 338 14 340 26
rect 348 14 350 26
rect 355 14 357 26
rect 365 14 367 26
rect 389 16 391 34
rect 402 6 404 27
rect 409 6 411 27
rect 430 6 432 34
rect 440 6 442 34
rect 450 6 452 34
rect 468 9 470 34
rect 475 9 477 34
rect 485 18 487 31
rect 498 6 500 31
rect 519 6 521 34
rect 529 6 531 34
rect 539 6 541 34
rect 557 9 559 34
rect 564 9 566 34
rect 574 18 576 31
rect 587 6 589 31
rect 607 26 609 34
rect 617 6 619 22
rect 624 6 626 22
rect 634 6 636 22
rect 641 6 643 22
rect 651 6 653 24
rect 671 16 673 34
<< polyct0 >>
rect 61 262 63 264
rect 36 247 38 249
rect 54 246 56 248
rect 107 255 109 257
rect 101 245 103 247
rect 157 252 159 254
rect 167 252 169 254
rect 196 255 198 257
rect 190 245 192 247
rect 246 252 248 254
rect 256 252 258 254
rect 295 252 297 254
rect 347 260 349 262
rect 322 244 324 246
rect 340 244 342 246
rect 440 261 442 263
rect 447 245 449 247
rect 512 261 514 263
rect 465 245 467 247
rect 487 245 489 247
rect 505 245 507 247
rect 576 261 578 263
rect 551 245 553 247
rect 569 245 571 247
rect 616 254 618 256
rect 657 253 659 255
rect 29 185 31 187
rect 70 184 72 186
rect 117 193 119 195
rect 135 193 137 195
rect 110 177 112 179
rect 181 193 183 195
rect 199 193 201 195
rect 221 193 223 195
rect 174 177 176 179
rect 239 193 241 195
rect 246 177 248 179
rect 346 194 348 196
rect 364 194 366 196
rect 339 178 341 180
rect 391 186 393 188
rect 430 186 432 188
rect 440 186 442 188
rect 496 193 498 195
rect 490 183 492 185
rect 519 186 521 188
rect 529 186 531 188
rect 585 193 587 195
rect 579 183 581 185
rect 632 192 634 194
rect 650 191 652 193
rect 625 176 627 178
rect 61 115 63 117
rect 36 100 38 102
rect 54 99 56 101
rect 107 108 109 110
rect 101 98 103 100
rect 157 105 159 107
rect 167 105 169 107
rect 196 108 198 110
rect 190 98 192 100
rect 246 105 248 107
rect 256 105 258 107
rect 295 105 297 107
rect 347 113 349 115
rect 322 97 324 99
rect 340 97 342 99
rect 440 114 442 116
rect 447 98 449 100
rect 512 114 514 116
rect 465 98 467 100
rect 487 98 489 100
rect 505 98 507 100
rect 576 114 578 116
rect 551 98 553 100
rect 569 98 571 100
rect 616 107 618 109
rect 657 106 659 108
rect 29 38 31 40
rect 70 37 72 39
rect 117 46 119 48
rect 135 46 137 48
rect 110 30 112 32
rect 181 46 183 48
rect 199 46 201 48
rect 221 46 223 48
rect 174 30 176 32
rect 239 46 241 48
rect 246 30 248 32
rect 346 47 348 49
rect 364 47 366 49
rect 339 31 341 33
rect 391 39 393 41
rect 430 39 432 41
rect 440 39 442 41
rect 496 46 498 48
rect 490 36 492 38
rect 519 39 521 41
rect 529 39 531 41
rect 585 46 587 48
rect 579 36 581 38
rect 632 45 634 47
rect 650 44 652 46
rect 625 29 627 31
<< polyct1 >>
rect 84 272 86 274
rect 13 252 15 254
rect 44 257 46 259
rect 71 252 73 254
rect 121 252 123 254
rect 140 252 142 254
rect 147 252 149 254
rect 275 259 277 261
rect 210 252 212 254
rect 229 252 231 254
rect 236 252 238 254
rect 370 270 372 272
rect 285 252 287 254
rect 330 254 332 256
rect 417 271 419 273
rect 393 260 395 262
rect 357 252 359 254
rect 535 271 537 273
rect 403 251 405 253
rect 430 253 432 255
rect 457 255 459 257
rect 495 255 497 257
rect 599 271 601 273
rect 522 253 524 255
rect 559 255 561 257
rect 667 277 669 279
rect 586 253 588 255
rect 626 261 628 263
rect 636 253 638 255
rect 676 245 678 247
rect 10 193 12 195
rect 50 185 52 187
rect 60 177 62 179
rect 100 185 102 187
rect 19 161 21 163
rect 127 183 129 185
rect 164 185 166 187
rect 87 167 89 169
rect 191 183 193 185
rect 229 183 231 185
rect 256 185 258 187
rect 283 187 285 189
rect 151 167 153 169
rect 329 186 331 188
rect 293 178 295 180
rect 269 167 271 169
rect 356 184 358 186
rect 401 186 403 188
rect 316 168 318 170
rect 450 186 452 188
rect 457 186 459 188
rect 476 186 478 188
rect 411 179 413 181
rect 539 186 541 188
rect 546 186 548 188
rect 565 186 567 188
rect 615 186 617 188
rect 642 181 644 183
rect 673 186 675 188
rect 602 166 604 168
rect 84 125 86 127
rect 13 105 15 107
rect 44 110 46 112
rect 71 105 73 107
rect 121 105 123 107
rect 140 105 142 107
rect 147 105 149 107
rect 275 112 277 114
rect 210 105 212 107
rect 229 105 231 107
rect 236 105 238 107
rect 370 123 372 125
rect 285 105 287 107
rect 330 107 332 109
rect 417 124 419 126
rect 393 113 395 115
rect 357 105 359 107
rect 535 124 537 126
rect 403 104 405 106
rect 430 106 432 108
rect 457 108 459 110
rect 495 108 497 110
rect 599 124 601 126
rect 522 106 524 108
rect 559 108 561 110
rect 667 130 669 132
rect 586 106 588 108
rect 626 114 628 116
rect 636 106 638 108
rect 676 98 678 100
rect 10 46 12 48
rect 50 38 52 40
rect 60 30 62 32
rect 100 38 102 40
rect 19 14 21 16
rect 127 36 129 38
rect 164 38 166 40
rect 87 20 89 22
rect 191 36 193 38
rect 229 36 231 38
rect 256 38 258 40
rect 283 40 285 42
rect 151 20 153 22
rect 329 39 331 41
rect 293 31 295 33
rect 269 20 271 22
rect 356 37 358 39
rect 401 39 403 41
rect 316 21 318 23
rect 450 39 452 41
rect 457 39 459 41
rect 476 39 478 41
rect 411 32 413 34
rect 539 39 541 41
rect 546 39 548 41
rect 565 39 567 41
rect 615 39 617 41
rect 642 34 644 36
rect 673 39 675 41
rect 602 19 604 21
<< ndifct0 >>
rect 6 240 8 242
rect 40 235 42 237
rect 57 235 59 237
rect 74 237 76 239
rect 84 237 86 239
rect 104 232 106 234
rect 114 235 116 237
rect 124 243 126 245
rect 134 243 136 245
rect 134 236 136 238
rect 144 236 146 238
rect 161 229 163 231
rect 193 232 195 234
rect 203 235 205 237
rect 213 243 215 245
rect 223 243 225 245
rect 223 236 225 238
rect 233 236 235 238
rect 282 243 284 245
rect 250 229 252 231
rect 386 242 388 244
rect 407 242 409 244
rect 272 230 274 232
rect 326 235 328 237
rect 343 235 345 237
rect 360 235 362 237
rect 370 235 372 237
rect 417 236 419 238
rect 427 236 429 238
rect 444 236 446 238
rect 461 236 463 238
rect 491 236 493 238
rect 508 236 510 238
rect 525 236 527 238
rect 535 236 537 238
rect 555 236 557 238
rect 572 236 574 238
rect 589 236 591 238
rect 599 236 601 238
rect 619 239 621 241
rect 629 239 631 241
rect 639 239 641 241
rect 291 230 293 232
rect 679 236 681 238
rect 7 202 9 204
rect 395 208 397 210
rect 47 199 49 201
rect 57 199 59 201
rect 67 199 69 201
rect 87 202 89 204
rect 97 202 99 204
rect 114 202 116 204
rect 131 202 133 204
rect 151 202 153 204
rect 161 202 163 204
rect 178 202 180 204
rect 195 202 197 204
rect 225 202 227 204
rect 242 202 244 204
rect 259 202 261 204
rect 269 202 271 204
rect 316 203 318 205
rect 326 203 328 205
rect 343 203 345 205
rect 360 203 362 205
rect 414 208 416 210
rect 279 196 281 198
rect 300 196 302 198
rect 436 209 438 211
rect 404 195 406 197
rect 453 202 455 204
rect 463 202 465 204
rect 463 195 465 197
rect 473 195 475 197
rect 483 203 485 205
rect 493 206 495 208
rect 525 209 527 211
rect 542 202 544 204
rect 552 202 554 204
rect 552 195 554 197
rect 562 195 564 197
rect 572 203 574 205
rect 582 206 584 208
rect 602 201 604 203
rect 612 201 614 203
rect 629 203 631 205
rect 646 203 648 205
rect 680 198 682 200
rect 6 93 8 95
rect 40 88 42 90
rect 57 88 59 90
rect 74 90 76 92
rect 84 90 86 92
rect 104 85 106 87
rect 114 88 116 90
rect 124 96 126 98
rect 134 96 136 98
rect 134 89 136 91
rect 144 89 146 91
rect 161 82 163 84
rect 193 85 195 87
rect 203 88 205 90
rect 213 96 215 98
rect 223 96 225 98
rect 223 89 225 91
rect 233 89 235 91
rect 282 96 284 98
rect 250 82 252 84
rect 386 95 388 97
rect 407 95 409 97
rect 272 83 274 85
rect 326 88 328 90
rect 343 88 345 90
rect 360 88 362 90
rect 370 88 372 90
rect 417 89 419 91
rect 427 89 429 91
rect 444 89 446 91
rect 461 89 463 91
rect 491 89 493 91
rect 508 89 510 91
rect 525 89 527 91
rect 535 89 537 91
rect 555 89 557 91
rect 572 89 574 91
rect 589 89 591 91
rect 599 89 601 91
rect 619 92 621 94
rect 629 92 631 94
rect 639 92 641 94
rect 291 83 293 85
rect 679 89 681 91
rect 7 55 9 57
rect 395 61 397 63
rect 47 52 49 54
rect 57 52 59 54
rect 67 52 69 54
rect 87 55 89 57
rect 97 55 99 57
rect 114 55 116 57
rect 131 55 133 57
rect 151 55 153 57
rect 161 55 163 57
rect 178 55 180 57
rect 195 55 197 57
rect 225 55 227 57
rect 242 55 244 57
rect 259 55 261 57
rect 269 55 271 57
rect 316 56 318 58
rect 326 56 328 58
rect 343 56 345 58
rect 360 56 362 58
rect 414 61 416 63
rect 279 49 281 51
rect 300 49 302 51
rect 436 62 438 64
rect 404 48 406 50
rect 453 55 455 57
rect 463 55 465 57
rect 463 48 465 50
rect 473 48 475 50
rect 483 56 485 58
rect 493 59 495 61
rect 525 62 527 64
rect 542 55 544 57
rect 552 55 554 57
rect 552 48 554 50
rect 562 48 564 50
rect 572 56 574 58
rect 582 59 584 61
rect 602 54 604 56
rect 612 54 614 56
rect 629 56 631 58
rect 646 56 648 58
rect 680 51 682 53
<< ndifct1 >>
rect 20 243 22 245
rect 30 238 32 240
rect 94 236 96 238
rect 172 236 174 238
rect 183 236 185 238
rect 261 236 263 238
rect 302 243 304 245
rect 397 242 399 244
rect 316 235 318 237
rect 471 236 473 238
rect 481 236 483 238
rect 545 236 547 238
rect 609 239 611 241
rect 650 239 652 241
rect 661 227 663 229
rect 25 211 27 213
rect 36 199 38 201
rect 77 199 79 201
rect 141 202 143 204
rect 205 202 207 204
rect 215 202 217 204
rect 370 203 372 205
rect 289 196 291 198
rect 384 195 386 197
rect 425 202 427 204
rect 503 202 505 204
rect 514 202 516 204
rect 592 202 594 204
rect 656 200 658 202
rect 666 195 668 197
rect 20 96 22 98
rect 30 91 32 93
rect 94 89 96 91
rect 172 89 174 91
rect 183 89 185 91
rect 261 89 263 91
rect 302 96 304 98
rect 397 95 399 97
rect 316 88 318 90
rect 471 89 473 91
rect 481 89 483 91
rect 545 89 547 91
rect 609 92 611 94
rect 650 92 652 94
rect 661 80 663 82
rect 25 64 27 66
rect 36 52 38 54
rect 77 52 79 54
rect 141 55 143 57
rect 205 55 207 57
rect 215 55 217 57
rect 370 56 372 58
rect 289 49 291 51
rect 384 48 386 50
rect 425 55 427 57
rect 503 55 505 57
rect 514 55 516 57
rect 592 55 594 57
rect 656 53 658 55
rect 666 48 668 50
<< ntiect1 >>
rect 7 286 9 288
rect 19 286 21 288
rect 301 286 303 288
rect 369 286 371 288
rect 418 287 420 289
rect 534 287 536 289
rect 598 287 600 289
rect 610 287 612 289
rect 651 287 653 289
rect 665 287 667 289
rect 679 287 681 289
rect 7 151 9 153
rect 21 151 23 153
rect 35 151 37 153
rect 76 151 78 153
rect 88 151 90 153
rect 152 151 154 153
rect 268 151 270 153
rect 317 152 319 154
rect 385 152 387 154
rect 667 152 669 154
rect 679 152 681 154
rect 7 139 9 141
rect 19 139 21 141
rect 301 139 303 141
rect 369 139 371 141
rect 418 140 420 142
rect 534 140 536 142
rect 598 140 600 142
rect 610 140 612 142
rect 651 140 653 142
rect 665 140 667 142
rect 679 140 681 142
rect 7 4 9 6
rect 21 4 23 6
rect 35 4 37 6
rect 76 4 78 6
rect 88 4 90 6
rect 152 4 154 6
rect 268 4 270 6
rect 317 5 319 7
rect 385 5 387 7
rect 667 5 669 7
rect 679 5 681 7
<< ptiect1 >>
rect 7 226 9 228
rect 19 226 21 228
rect 301 226 303 228
rect 387 226 389 228
rect 407 226 409 228
rect 610 227 612 229
rect 638 227 640 229
rect 651 227 653 229
rect 35 211 37 213
rect 48 211 50 213
rect 76 211 78 213
rect 279 212 281 214
rect 299 212 301 214
rect 385 212 387 214
rect 667 212 669 214
rect 679 212 681 214
rect 7 79 9 81
rect 19 79 21 81
rect 301 79 303 81
rect 387 79 389 81
rect 407 79 409 81
rect 610 80 612 82
rect 638 80 640 82
rect 651 80 653 82
rect 35 64 37 66
rect 48 64 50 66
rect 76 64 78 66
rect 279 65 281 67
rect 299 65 301 67
rect 385 65 387 67
rect 667 65 669 67
rect 679 65 681 67
<< pdifct0 >>
rect 9 276 11 278
rect 40 283 42 285
rect 57 273 59 275
rect 74 283 76 285
rect 84 261 86 263
rect 105 283 107 285
rect 117 264 119 266
rect 140 283 142 285
rect 140 276 142 278
rect 152 275 154 277
rect 152 268 154 270
rect 162 283 164 285
rect 162 276 164 278
rect 194 283 196 285
rect 206 264 208 266
rect 229 283 231 285
rect 229 276 231 278
rect 241 275 243 277
rect 241 268 243 270
rect 251 283 253 285
rect 251 276 253 278
rect 272 276 274 278
rect 291 283 293 285
rect 326 275 328 277
rect 343 269 345 271
rect 360 275 362 277
rect 408 283 410 285
rect 621 284 623 286
rect 408 276 410 278
rect 427 276 429 278
rect 370 261 372 263
rect 444 270 446 272
rect 461 276 463 278
rect 491 276 493 278
rect 508 270 510 272
rect 525 276 527 278
rect 417 262 419 264
rect 555 276 557 278
rect 572 270 574 272
rect 589 276 591 278
rect 535 262 537 264
rect 639 277 641 279
rect 599 262 601 264
rect 660 262 662 264
rect 670 262 672 264
rect 680 266 682 268
rect 6 172 8 174
rect 16 176 18 178
rect 26 176 28 178
rect 87 176 89 178
rect 47 161 49 163
rect 151 176 153 178
rect 97 162 99 164
rect 114 168 116 170
rect 131 162 133 164
rect 269 176 271 178
rect 161 162 163 164
rect 178 168 180 170
rect 195 162 197 164
rect 225 162 227 164
rect 242 168 244 170
rect 316 177 318 179
rect 259 162 261 164
rect 278 162 280 164
rect 65 154 67 156
rect 278 155 280 157
rect 326 163 328 165
rect 343 169 345 171
rect 360 163 362 165
rect 395 155 397 157
rect 414 162 416 164
rect 435 162 437 164
rect 435 155 437 157
rect 445 170 447 172
rect 445 163 447 165
rect 457 162 459 164
rect 457 155 459 157
rect 480 174 482 176
rect 492 155 494 157
rect 524 162 526 164
rect 524 155 526 157
rect 534 170 536 172
rect 534 163 536 165
rect 546 162 548 164
rect 546 155 548 157
rect 569 174 571 176
rect 581 155 583 157
rect 602 177 604 179
rect 612 155 614 157
rect 629 165 631 167
rect 646 155 648 157
rect 677 162 679 164
rect 9 129 11 131
rect 40 136 42 138
rect 57 126 59 128
rect 74 136 76 138
rect 84 114 86 116
rect 105 136 107 138
rect 117 117 119 119
rect 140 136 142 138
rect 140 129 142 131
rect 152 128 154 130
rect 152 121 154 123
rect 162 136 164 138
rect 162 129 164 131
rect 194 136 196 138
rect 206 117 208 119
rect 229 136 231 138
rect 229 129 231 131
rect 241 128 243 130
rect 241 121 243 123
rect 251 136 253 138
rect 251 129 253 131
rect 272 129 274 131
rect 291 136 293 138
rect 326 128 328 130
rect 343 122 345 124
rect 360 128 362 130
rect 408 136 410 138
rect 621 137 623 139
rect 408 129 410 131
rect 427 129 429 131
rect 370 114 372 116
rect 444 123 446 125
rect 461 129 463 131
rect 491 129 493 131
rect 508 123 510 125
rect 525 129 527 131
rect 417 115 419 117
rect 555 129 557 131
rect 572 123 574 125
rect 589 129 591 131
rect 535 115 537 117
rect 639 130 641 132
rect 599 115 601 117
rect 660 115 662 117
rect 670 115 672 117
rect 680 119 682 121
rect 6 25 8 27
rect 16 29 18 31
rect 26 29 28 31
rect 87 29 89 31
rect 47 14 49 16
rect 151 29 153 31
rect 97 15 99 17
rect 114 21 116 23
rect 131 15 133 17
rect 269 29 271 31
rect 161 15 163 17
rect 178 21 180 23
rect 195 15 197 17
rect 225 15 227 17
rect 242 21 244 23
rect 316 30 318 32
rect 259 15 261 17
rect 278 15 280 17
rect 65 7 67 9
rect 278 8 280 10
rect 326 16 328 18
rect 343 22 345 24
rect 360 16 362 18
rect 395 8 397 10
rect 414 15 416 17
rect 435 15 437 17
rect 435 8 437 10
rect 445 23 447 25
rect 445 16 447 18
rect 457 15 459 17
rect 457 8 459 10
rect 480 27 482 29
rect 492 8 494 10
rect 524 15 526 17
rect 524 8 526 10
rect 534 23 536 25
rect 534 16 536 18
rect 546 15 548 17
rect 546 8 548 10
rect 569 27 571 29
rect 581 8 583 10
rect 602 30 604 32
rect 612 8 614 10
rect 629 18 631 20
rect 646 8 648 10
rect 677 15 679 17
<< pdifct1 >>
rect 30 276 32 278
rect 20 268 22 270
rect 20 261 22 263
rect 94 271 96 273
rect 94 264 96 266
rect 172 268 174 270
rect 172 261 174 263
rect 183 271 185 273
rect 183 264 185 266
rect 261 268 263 270
rect 261 261 263 263
rect 302 273 304 275
rect 302 266 304 268
rect 316 269 318 271
rect 389 277 391 279
rect 471 270 473 272
rect 481 270 483 272
rect 545 270 547 272
rect 609 275 611 277
rect 650 262 652 264
rect 36 176 38 178
rect 77 163 79 165
rect 141 168 143 170
rect 205 168 207 170
rect 215 168 217 170
rect 297 161 299 163
rect 370 169 372 171
rect 384 172 386 174
rect 384 165 386 167
rect 425 177 427 179
rect 425 170 427 172
rect 503 174 505 176
rect 503 167 505 169
rect 514 177 516 179
rect 514 170 516 172
rect 592 174 594 176
rect 592 167 594 169
rect 666 177 668 179
rect 666 170 668 172
rect 656 162 658 164
rect 30 129 32 131
rect 20 121 22 123
rect 20 114 22 116
rect 94 124 96 126
rect 94 117 96 119
rect 172 121 174 123
rect 172 114 174 116
rect 183 124 185 126
rect 183 117 185 119
rect 261 121 263 123
rect 261 114 263 116
rect 302 126 304 128
rect 302 119 304 121
rect 316 122 318 124
rect 389 130 391 132
rect 471 123 473 125
rect 481 123 483 125
rect 545 123 547 125
rect 609 128 611 130
rect 650 115 652 117
rect 36 29 38 31
rect 77 16 79 18
rect 141 21 143 23
rect 205 21 207 23
rect 215 21 217 23
rect 297 14 299 16
rect 370 22 372 24
rect 384 25 386 27
rect 384 18 386 20
rect 425 30 427 32
rect 425 23 427 25
rect 503 27 505 29
rect 503 20 505 22
rect 514 30 516 32
rect 514 23 516 25
rect 592 27 594 29
rect 592 20 594 22
rect 666 30 668 32
rect 666 23 668 25
rect 656 15 658 17
<< alu0 >>
rect 7 278 13 285
rect 38 283 40 285
rect 42 283 44 285
rect 38 282 44 283
rect 73 283 74 285
rect 76 283 77 285
rect 73 281 77 283
rect 103 283 105 285
rect 107 283 109 285
rect 103 282 109 283
rect 138 283 140 285
rect 142 283 144 285
rect 7 276 9 278
rect 11 276 13 278
rect 7 275 13 276
rect 48 275 61 276
rect 19 259 20 266
rect 5 242 9 244
rect 5 240 6 242
rect 8 240 9 242
rect 19 241 20 247
rect 5 229 9 240
rect 48 273 57 275
rect 59 273 61 275
rect 48 272 61 273
rect 36 268 52 272
rect 36 251 40 268
rect 138 278 144 283
rect 160 283 162 285
rect 164 283 166 285
rect 138 276 140 278
rect 142 276 144 278
rect 138 275 144 276
rect 151 277 155 279
rect 151 275 152 277
rect 154 275 155 277
rect 160 278 166 283
rect 192 283 194 285
rect 196 283 198 285
rect 192 282 198 283
rect 227 283 229 285
rect 231 283 233 285
rect 160 276 162 278
rect 164 276 166 278
rect 160 275 166 276
rect 227 278 233 283
rect 249 283 251 285
rect 253 283 255 285
rect 227 276 229 278
rect 231 276 233 278
rect 227 275 233 276
rect 240 277 244 279
rect 240 275 241 277
rect 243 275 244 277
rect 249 278 255 283
rect 289 283 291 285
rect 293 283 295 285
rect 289 282 295 283
rect 249 276 251 278
rect 253 276 255 278
rect 249 275 255 276
rect 270 278 287 279
rect 270 276 272 278
rect 274 276 287 278
rect 270 275 287 276
rect 108 271 132 275
rect 151 271 155 275
rect 60 264 64 266
rect 43 255 44 261
rect 60 262 61 264
rect 63 263 88 264
rect 63 262 84 263
rect 60 261 84 262
rect 86 261 88 263
rect 60 260 88 261
rect 35 249 40 251
rect 60 250 64 260
rect 35 247 36 249
rect 38 247 40 249
rect 53 248 64 250
rect 35 245 50 247
rect 36 243 50 245
rect 53 246 54 248
rect 56 246 64 248
rect 53 244 64 246
rect 39 237 43 239
rect 39 235 40 237
rect 42 235 43 237
rect 39 229 43 235
rect 46 238 50 243
rect 84 240 88 260
rect 72 239 78 240
rect 46 237 61 238
rect 46 235 57 237
rect 59 235 61 237
rect 46 234 61 235
rect 72 237 74 239
rect 76 237 78 239
rect 72 229 78 237
rect 82 239 88 240
rect 82 237 84 239
rect 86 237 88 239
rect 82 236 88 237
rect 106 267 112 271
rect 128 270 168 271
rect 128 268 152 270
rect 154 268 168 270
rect 106 257 110 267
rect 116 266 120 268
rect 128 267 168 268
rect 116 264 117 266
rect 119 264 120 266
rect 116 263 120 264
rect 106 255 107 257
rect 109 255 110 257
rect 106 253 110 255
rect 113 259 120 263
rect 113 248 117 259
rect 156 254 160 259
rect 156 252 157 254
rect 159 252 160 254
rect 99 247 117 248
rect 99 245 101 247
rect 103 246 117 247
rect 103 245 128 246
rect 99 244 124 245
rect 113 243 124 244
rect 126 243 128 245
rect 113 242 128 243
rect 133 245 137 247
rect 133 243 134 245
rect 136 243 137 245
rect 133 238 137 243
rect 156 250 160 252
rect 164 256 168 267
rect 164 254 170 256
rect 164 252 167 254
rect 169 252 170 254
rect 164 250 170 252
rect 164 247 168 250
rect 148 243 168 247
rect 148 239 152 243
rect 112 237 134 238
rect 103 234 107 236
rect 112 235 114 237
rect 116 236 134 237
rect 136 236 137 238
rect 116 235 137 236
rect 142 238 152 239
rect 142 236 144 238
rect 146 236 152 238
rect 142 235 152 236
rect 197 271 221 275
rect 240 271 244 275
rect 195 267 201 271
rect 217 270 257 271
rect 217 268 241 270
rect 243 268 257 270
rect 195 257 199 267
rect 205 266 209 268
rect 217 267 257 268
rect 205 264 206 266
rect 208 264 209 266
rect 205 263 209 264
rect 195 255 196 257
rect 198 255 199 257
rect 195 253 199 255
rect 202 259 209 263
rect 202 248 206 259
rect 245 254 249 259
rect 245 252 246 254
rect 248 252 249 254
rect 188 247 206 248
rect 188 245 190 247
rect 192 246 206 247
rect 192 245 217 246
rect 188 244 213 245
rect 202 243 213 244
rect 215 243 217 245
rect 202 242 217 243
rect 222 245 226 247
rect 222 243 223 245
rect 225 243 226 245
rect 222 238 226 243
rect 245 250 249 252
rect 253 256 257 267
rect 283 271 287 275
rect 283 267 298 271
rect 253 254 259 256
rect 253 252 256 254
rect 258 252 259 254
rect 253 250 259 252
rect 253 247 257 250
rect 237 243 257 247
rect 237 239 241 243
rect 273 258 279 259
rect 294 254 298 267
rect 301 264 302 275
rect 324 277 330 285
rect 324 275 326 277
rect 328 275 330 277
rect 324 274 330 275
rect 358 277 364 285
rect 407 283 408 285
rect 410 283 411 285
rect 358 275 360 277
rect 362 275 364 277
rect 358 274 364 275
rect 294 252 295 254
rect 297 252 298 254
rect 294 246 298 252
rect 280 245 298 246
rect 280 243 282 245
rect 284 243 298 245
rect 280 242 298 243
rect 341 271 347 272
rect 330 269 343 271
rect 345 269 347 271
rect 330 267 347 269
rect 407 278 411 283
rect 407 276 408 278
rect 410 276 411 278
rect 201 237 223 238
rect 112 234 137 235
rect 192 234 196 236
rect 201 235 203 237
rect 205 236 223 237
rect 225 236 226 238
rect 205 235 226 236
rect 231 238 241 239
rect 231 236 233 238
rect 235 236 241 238
rect 231 235 241 236
rect 330 264 334 267
rect 321 260 334 264
rect 346 263 374 264
rect 321 246 325 260
rect 346 262 370 263
rect 346 260 347 262
rect 349 261 370 262
rect 372 261 374 263
rect 349 260 374 261
rect 346 248 350 260
rect 339 246 350 248
rect 321 244 322 246
rect 324 244 336 246
rect 321 242 336 244
rect 339 244 340 246
rect 342 244 350 246
rect 339 242 350 244
rect 201 234 226 235
rect 325 237 329 239
rect 325 235 326 237
rect 328 235 329 237
rect 103 232 104 234
rect 106 232 107 234
rect 192 232 193 234
rect 195 232 196 234
rect 270 232 276 233
rect 103 229 107 232
rect 159 231 165 232
rect 159 229 161 231
rect 163 229 165 231
rect 192 229 196 232
rect 248 231 254 232
rect 248 229 250 231
rect 252 229 254 231
rect 270 230 272 232
rect 274 230 276 232
rect 270 229 276 230
rect 289 232 295 233
rect 289 230 291 232
rect 293 230 295 232
rect 289 229 295 230
rect 325 229 329 235
rect 332 238 336 242
rect 370 238 374 260
rect 407 274 411 276
rect 425 278 431 286
rect 425 276 427 278
rect 429 276 431 278
rect 425 275 431 276
rect 459 278 465 286
rect 459 276 461 278
rect 463 276 465 278
rect 459 275 465 276
rect 489 278 495 286
rect 489 276 491 278
rect 493 276 495 278
rect 489 275 495 276
rect 523 278 529 286
rect 523 276 525 278
rect 527 276 529 278
rect 523 275 529 276
rect 553 278 559 286
rect 553 276 555 278
rect 557 276 559 278
rect 553 275 559 276
rect 587 278 593 286
rect 619 284 621 286
rect 623 284 625 286
rect 619 283 625 284
rect 587 276 589 278
rect 591 276 593 278
rect 587 275 593 276
rect 442 272 448 273
rect 442 270 444 272
rect 446 270 459 272
rect 442 268 459 270
rect 455 265 459 268
rect 415 264 443 265
rect 415 262 417 264
rect 419 263 443 264
rect 419 262 440 263
rect 415 261 440 262
rect 442 261 443 263
rect 332 237 347 238
rect 332 235 343 237
rect 345 235 347 237
rect 332 234 347 235
rect 358 237 364 238
rect 358 235 360 237
rect 362 235 364 237
rect 358 229 364 235
rect 368 237 374 238
rect 368 235 370 237
rect 372 235 374 237
rect 368 234 374 235
rect 385 244 389 246
rect 385 242 386 244
rect 388 242 389 244
rect 385 230 389 242
rect 406 244 411 246
rect 406 242 407 244
rect 409 242 411 244
rect 406 240 411 242
rect 407 230 411 240
rect 415 239 419 261
rect 439 249 443 261
rect 455 261 468 265
rect 439 247 450 249
rect 464 247 468 261
rect 439 245 447 247
rect 449 245 450 247
rect 439 243 450 245
rect 453 245 465 247
rect 467 245 468 247
rect 453 243 468 245
rect 453 239 457 243
rect 415 238 421 239
rect 415 236 417 238
rect 419 236 421 238
rect 415 235 421 236
rect 425 238 431 239
rect 425 236 427 238
rect 429 236 431 238
rect 425 230 431 236
rect 442 238 457 239
rect 442 236 444 238
rect 446 236 457 238
rect 442 235 457 236
rect 460 238 464 240
rect 460 236 461 238
rect 463 236 464 238
rect 460 230 464 236
rect 506 272 512 273
rect 495 270 508 272
rect 510 270 512 272
rect 495 268 512 270
rect 570 272 576 273
rect 559 270 572 272
rect 574 270 576 272
rect 559 268 576 270
rect 623 279 643 280
rect 623 277 639 279
rect 641 277 643 279
rect 623 276 643 277
rect 495 265 499 268
rect 486 261 499 265
rect 511 264 539 265
rect 486 247 490 261
rect 511 263 535 264
rect 511 261 512 263
rect 514 262 535 263
rect 537 262 539 264
rect 514 261 539 262
rect 511 249 515 261
rect 504 247 515 249
rect 486 245 487 247
rect 489 245 501 247
rect 486 243 501 245
rect 504 245 505 247
rect 507 245 515 247
rect 504 243 515 245
rect 490 238 494 240
rect 490 236 491 238
rect 493 236 494 238
rect 490 230 494 236
rect 497 239 501 243
rect 535 239 539 261
rect 497 238 512 239
rect 497 236 508 238
rect 510 236 512 238
rect 497 235 512 236
rect 523 238 529 239
rect 523 236 525 238
rect 527 236 529 238
rect 523 230 529 236
rect 533 238 539 239
rect 533 236 535 238
rect 537 236 539 238
rect 533 235 539 236
rect 559 265 563 268
rect 550 261 563 265
rect 575 264 603 265
rect 550 247 554 261
rect 575 263 599 264
rect 575 261 576 263
rect 578 262 599 263
rect 601 262 603 264
rect 578 261 603 262
rect 575 249 579 261
rect 568 247 579 249
rect 550 245 551 247
rect 553 245 565 247
rect 550 243 565 245
rect 568 245 569 247
rect 571 245 579 247
rect 568 243 579 245
rect 554 238 558 240
rect 554 236 555 238
rect 557 236 558 238
rect 554 230 558 236
rect 561 239 565 243
rect 599 239 603 261
rect 561 238 576 239
rect 561 236 572 238
rect 574 236 576 238
rect 561 235 576 236
rect 587 238 593 239
rect 587 236 589 238
rect 591 236 593 238
rect 587 230 593 236
rect 597 238 603 239
rect 597 236 599 238
rect 601 236 603 238
rect 597 235 603 236
rect 611 273 612 276
rect 623 272 627 276
rect 615 268 627 272
rect 615 256 619 268
rect 615 254 616 256
rect 618 254 619 256
rect 615 249 619 254
rect 615 245 632 249
rect 617 241 623 242
rect 617 239 619 241
rect 621 239 623 241
rect 617 230 623 239
rect 628 241 632 245
rect 652 260 653 266
rect 656 265 660 286
rect 679 281 683 286
rect 679 268 683 277
rect 679 266 680 268
rect 682 266 683 268
rect 656 264 664 265
rect 656 262 660 264
rect 662 262 664 264
rect 656 261 664 262
rect 668 264 674 265
rect 679 264 683 266
rect 668 262 670 264
rect 672 262 674 264
rect 668 256 674 262
rect 655 255 674 256
rect 655 253 657 255
rect 659 253 674 255
rect 655 252 674 253
rect 628 239 629 241
rect 631 239 632 241
rect 628 237 632 239
rect 637 241 643 242
rect 637 239 639 241
rect 641 239 643 241
rect 637 230 643 239
rect 652 241 653 243
rect 664 239 668 252
rect 664 238 683 239
rect 664 236 679 238
rect 681 236 683 238
rect 664 235 683 236
rect 5 204 24 205
rect 5 202 7 204
rect 9 202 24 204
rect 5 201 24 202
rect 20 188 24 201
rect 35 197 36 199
rect 45 201 51 210
rect 45 199 47 201
rect 49 199 51 201
rect 45 198 51 199
rect 56 201 60 203
rect 56 199 57 201
rect 59 199 60 201
rect 14 187 33 188
rect 14 185 29 187
rect 31 185 33 187
rect 14 184 33 185
rect 14 178 20 184
rect 14 176 16 178
rect 18 176 20 178
rect 5 174 9 176
rect 14 175 20 176
rect 24 178 32 179
rect 24 176 26 178
rect 28 176 32 178
rect 24 175 32 176
rect 5 172 6 174
rect 8 172 9 174
rect 5 154 9 172
rect 28 154 32 175
rect 35 174 36 180
rect 56 195 60 199
rect 65 201 71 210
rect 65 199 67 201
rect 69 199 71 201
rect 65 198 71 199
rect 56 191 73 195
rect 69 186 73 191
rect 69 184 70 186
rect 72 184 73 186
rect 69 172 73 184
rect 61 168 73 172
rect 61 164 65 168
rect 76 164 77 167
rect 85 204 91 205
rect 85 202 87 204
rect 89 202 91 204
rect 85 201 91 202
rect 95 204 101 210
rect 95 202 97 204
rect 99 202 101 204
rect 95 201 101 202
rect 112 204 127 205
rect 112 202 114 204
rect 116 202 127 204
rect 112 201 127 202
rect 85 179 89 201
rect 123 197 127 201
rect 130 204 134 210
rect 130 202 131 204
rect 133 202 134 204
rect 130 200 134 202
rect 109 195 120 197
rect 109 193 117 195
rect 119 193 120 195
rect 123 195 138 197
rect 123 193 135 195
rect 137 193 138 195
rect 109 191 120 193
rect 109 179 113 191
rect 85 178 110 179
rect 85 176 87 178
rect 89 177 110 178
rect 112 177 113 179
rect 89 176 113 177
rect 134 179 138 193
rect 85 175 113 176
rect 125 175 138 179
rect 125 172 129 175
rect 149 204 155 205
rect 149 202 151 204
rect 153 202 155 204
rect 149 201 155 202
rect 159 204 165 210
rect 159 202 161 204
rect 163 202 165 204
rect 159 201 165 202
rect 176 204 191 205
rect 176 202 178 204
rect 180 202 191 204
rect 176 201 191 202
rect 149 179 153 201
rect 187 197 191 201
rect 194 204 198 210
rect 194 202 195 204
rect 197 202 198 204
rect 194 200 198 202
rect 173 195 184 197
rect 173 193 181 195
rect 183 193 184 195
rect 187 195 202 197
rect 187 193 199 195
rect 201 193 202 195
rect 173 191 184 193
rect 173 179 177 191
rect 149 178 174 179
rect 149 176 151 178
rect 153 177 174 178
rect 176 177 177 179
rect 153 176 177 177
rect 198 179 202 193
rect 149 175 177 176
rect 189 175 202 179
rect 189 172 193 175
rect 45 163 65 164
rect 45 161 47 163
rect 49 161 65 163
rect 45 160 65 161
rect 112 170 129 172
rect 112 168 114 170
rect 116 168 129 170
rect 112 167 118 168
rect 176 170 193 172
rect 176 168 178 170
rect 180 168 193 170
rect 176 167 182 168
rect 224 204 228 210
rect 224 202 225 204
rect 227 202 228 204
rect 224 200 228 202
rect 231 204 246 205
rect 231 202 242 204
rect 244 202 246 204
rect 231 201 246 202
rect 257 204 263 210
rect 257 202 259 204
rect 261 202 263 204
rect 257 201 263 202
rect 267 204 273 205
rect 267 202 269 204
rect 271 202 273 204
rect 267 201 273 202
rect 231 197 235 201
rect 220 195 235 197
rect 220 193 221 195
rect 223 193 235 195
rect 238 195 249 197
rect 238 193 239 195
rect 241 193 249 195
rect 220 179 224 193
rect 238 191 249 193
rect 220 175 233 179
rect 245 179 249 191
rect 269 179 273 201
rect 277 200 281 210
rect 277 198 282 200
rect 277 196 279 198
rect 281 196 282 198
rect 277 194 282 196
rect 299 198 303 210
rect 299 196 300 198
rect 302 196 303 198
rect 299 194 303 196
rect 314 205 320 206
rect 314 203 316 205
rect 318 203 320 205
rect 314 202 320 203
rect 324 205 330 211
rect 324 203 326 205
rect 328 203 330 205
rect 324 202 330 203
rect 341 205 356 206
rect 341 203 343 205
rect 345 203 356 205
rect 341 202 356 203
rect 245 177 246 179
rect 248 178 273 179
rect 248 177 269 178
rect 245 176 269 177
rect 271 176 273 178
rect 245 175 273 176
rect 229 172 233 175
rect 229 170 246 172
rect 229 168 242 170
rect 244 168 246 170
rect 240 167 246 168
rect 95 164 101 165
rect 95 162 97 164
rect 99 162 101 164
rect 63 156 69 157
rect 63 154 65 156
rect 67 154 69 156
rect 95 154 101 162
rect 129 164 135 165
rect 129 162 131 164
rect 133 162 135 164
rect 129 154 135 162
rect 159 164 165 165
rect 159 162 161 164
rect 163 162 165 164
rect 159 154 165 162
rect 193 164 199 165
rect 193 162 195 164
rect 197 162 199 164
rect 193 154 199 162
rect 223 164 229 165
rect 223 162 225 164
rect 227 162 229 164
rect 223 154 229 162
rect 257 164 263 165
rect 257 162 259 164
rect 261 162 263 164
rect 257 154 263 162
rect 277 164 281 166
rect 314 180 318 202
rect 352 198 356 202
rect 359 205 363 211
rect 393 210 399 211
rect 393 208 395 210
rect 397 208 399 210
rect 393 207 399 208
rect 412 210 418 211
rect 412 208 414 210
rect 416 208 418 210
rect 434 209 436 211
rect 438 209 440 211
rect 434 208 440 209
rect 492 208 496 211
rect 523 209 525 211
rect 527 209 529 211
rect 523 208 529 209
rect 581 208 585 211
rect 412 207 418 208
rect 492 206 493 208
rect 495 206 496 208
rect 581 206 582 208
rect 584 206 585 208
rect 359 203 360 205
rect 362 203 363 205
rect 359 201 363 203
rect 462 205 487 206
rect 338 196 349 198
rect 338 194 346 196
rect 348 194 349 196
rect 352 196 367 198
rect 352 194 364 196
rect 366 194 367 196
rect 338 192 349 194
rect 338 180 342 192
rect 314 179 339 180
rect 314 177 316 179
rect 318 178 339 179
rect 341 178 342 180
rect 318 177 342 178
rect 363 180 367 194
rect 314 176 342 177
rect 354 176 367 180
rect 447 204 457 205
rect 447 202 453 204
rect 455 202 457 204
rect 447 201 457 202
rect 462 204 483 205
rect 462 202 463 204
rect 465 203 483 204
rect 485 203 487 205
rect 492 204 496 206
rect 551 205 576 206
rect 465 202 487 203
rect 354 173 358 176
rect 277 162 278 164
rect 280 162 281 164
rect 277 157 281 162
rect 341 171 358 173
rect 341 169 343 171
rect 345 169 358 171
rect 341 168 347 169
rect 390 197 408 198
rect 390 195 404 197
rect 406 195 408 197
rect 390 194 408 195
rect 390 188 394 194
rect 390 186 391 188
rect 393 186 394 188
rect 324 165 330 166
rect 324 163 326 165
rect 328 163 330 165
rect 277 155 278 157
rect 280 155 281 157
rect 324 155 330 163
rect 358 165 364 166
rect 358 163 360 165
rect 362 163 364 165
rect 358 155 364 163
rect 386 165 387 176
rect 390 173 394 186
rect 409 181 415 182
rect 447 197 451 201
rect 431 193 451 197
rect 431 190 435 193
rect 429 188 435 190
rect 429 186 430 188
rect 432 186 435 188
rect 429 184 435 186
rect 390 169 405 173
rect 401 165 405 169
rect 431 173 435 184
rect 439 188 443 190
rect 462 197 466 202
rect 462 195 463 197
rect 465 195 466 197
rect 462 193 466 195
rect 471 197 486 198
rect 471 195 473 197
rect 475 196 486 197
rect 475 195 500 196
rect 471 194 496 195
rect 482 193 496 194
rect 498 193 500 195
rect 482 192 500 193
rect 439 186 440 188
rect 442 186 443 188
rect 439 181 443 186
rect 482 181 486 192
rect 479 177 486 181
rect 489 185 493 187
rect 489 183 490 185
rect 492 183 493 185
rect 479 176 483 177
rect 479 174 480 176
rect 482 174 483 176
rect 431 172 471 173
rect 479 172 483 174
rect 489 173 493 183
rect 431 170 445 172
rect 447 170 471 172
rect 431 169 471 170
rect 487 169 493 173
rect 444 165 448 169
rect 467 165 491 169
rect 536 204 546 205
rect 536 202 542 204
rect 544 202 546 204
rect 536 201 546 202
rect 551 204 572 205
rect 551 202 552 204
rect 554 203 572 204
rect 574 203 576 205
rect 581 204 585 206
rect 554 202 576 203
rect 536 197 540 201
rect 520 193 540 197
rect 520 190 524 193
rect 518 188 524 190
rect 518 186 519 188
rect 521 186 524 188
rect 518 184 524 186
rect 520 173 524 184
rect 528 188 532 190
rect 551 197 555 202
rect 551 195 552 197
rect 554 195 555 197
rect 551 193 555 195
rect 560 197 575 198
rect 560 195 562 197
rect 564 196 575 197
rect 564 195 589 196
rect 560 194 585 195
rect 571 193 585 194
rect 587 193 589 195
rect 571 192 589 193
rect 528 186 529 188
rect 531 186 532 188
rect 528 181 532 186
rect 571 181 575 192
rect 568 177 575 181
rect 578 185 582 187
rect 578 183 579 185
rect 581 183 582 185
rect 568 176 572 177
rect 568 174 569 176
rect 571 174 572 176
rect 520 172 560 173
rect 568 172 572 174
rect 578 173 582 183
rect 520 170 534 172
rect 536 170 560 172
rect 520 169 560 170
rect 576 169 582 173
rect 600 203 606 204
rect 600 201 602 203
rect 604 201 606 203
rect 600 200 606 201
rect 610 203 616 211
rect 610 201 612 203
rect 614 201 616 203
rect 627 205 642 206
rect 627 203 629 205
rect 631 203 642 205
rect 627 202 642 203
rect 610 200 616 201
rect 600 180 604 200
rect 638 197 642 202
rect 645 205 649 211
rect 645 203 646 205
rect 648 203 649 205
rect 645 201 649 203
rect 624 194 635 196
rect 624 192 632 194
rect 634 192 635 194
rect 638 195 652 197
rect 638 193 653 195
rect 624 190 635 192
rect 648 191 650 193
rect 652 191 653 193
rect 624 180 628 190
rect 648 189 653 191
rect 600 179 628 180
rect 600 177 602 179
rect 604 178 628 179
rect 604 177 625 178
rect 600 176 625 177
rect 627 176 628 178
rect 644 179 645 185
rect 624 174 628 176
rect 533 165 537 169
rect 556 165 580 169
rect 401 164 418 165
rect 401 162 414 164
rect 416 162 418 164
rect 401 161 418 162
rect 433 164 439 165
rect 433 162 435 164
rect 437 162 439 164
rect 393 157 399 158
rect 393 155 395 157
rect 397 155 399 157
rect 433 157 439 162
rect 444 163 445 165
rect 447 163 448 165
rect 444 161 448 163
rect 455 164 461 165
rect 455 162 457 164
rect 459 162 461 164
rect 433 155 435 157
rect 437 155 439 157
rect 455 157 461 162
rect 522 164 528 165
rect 522 162 524 164
rect 526 162 528 164
rect 455 155 457 157
rect 459 155 461 157
rect 490 157 496 158
rect 490 155 492 157
rect 494 155 496 157
rect 522 157 528 162
rect 533 163 534 165
rect 536 163 537 165
rect 533 161 537 163
rect 544 164 550 165
rect 544 162 546 164
rect 548 162 550 164
rect 522 155 524 157
rect 526 155 528 157
rect 544 157 550 162
rect 648 172 652 189
rect 636 168 652 172
rect 627 167 640 168
rect 627 165 629 167
rect 631 165 640 167
rect 679 200 683 211
rect 668 193 669 199
rect 679 198 680 200
rect 682 198 683 200
rect 679 196 683 198
rect 668 174 669 181
rect 627 164 640 165
rect 675 164 681 165
rect 675 162 677 164
rect 679 162 681 164
rect 544 155 546 157
rect 548 155 550 157
rect 579 157 585 158
rect 579 155 581 157
rect 583 155 585 157
rect 611 157 615 159
rect 611 155 612 157
rect 614 155 615 157
rect 644 157 650 158
rect 644 155 646 157
rect 648 155 650 157
rect 675 155 681 162
rect 7 131 13 138
rect 38 136 40 138
rect 42 136 44 138
rect 38 135 44 136
rect 73 136 74 138
rect 76 136 77 138
rect 73 134 77 136
rect 103 136 105 138
rect 107 136 109 138
rect 103 135 109 136
rect 138 136 140 138
rect 142 136 144 138
rect 7 129 9 131
rect 11 129 13 131
rect 7 128 13 129
rect 48 128 61 129
rect 19 112 20 119
rect 5 95 9 97
rect 5 93 6 95
rect 8 93 9 95
rect 19 94 20 100
rect 5 82 9 93
rect 48 126 57 128
rect 59 126 61 128
rect 48 125 61 126
rect 36 121 52 125
rect 36 104 40 121
rect 138 131 144 136
rect 160 136 162 138
rect 164 136 166 138
rect 138 129 140 131
rect 142 129 144 131
rect 138 128 144 129
rect 151 130 155 132
rect 151 128 152 130
rect 154 128 155 130
rect 160 131 166 136
rect 192 136 194 138
rect 196 136 198 138
rect 192 135 198 136
rect 227 136 229 138
rect 231 136 233 138
rect 160 129 162 131
rect 164 129 166 131
rect 160 128 166 129
rect 227 131 233 136
rect 249 136 251 138
rect 253 136 255 138
rect 227 129 229 131
rect 231 129 233 131
rect 227 128 233 129
rect 240 130 244 132
rect 240 128 241 130
rect 243 128 244 130
rect 249 131 255 136
rect 289 136 291 138
rect 293 136 295 138
rect 289 135 295 136
rect 249 129 251 131
rect 253 129 255 131
rect 249 128 255 129
rect 270 131 287 132
rect 270 129 272 131
rect 274 129 287 131
rect 270 128 287 129
rect 108 124 132 128
rect 151 124 155 128
rect 60 117 64 119
rect 43 108 44 114
rect 60 115 61 117
rect 63 116 88 117
rect 63 115 84 116
rect 60 114 84 115
rect 86 114 88 116
rect 60 113 88 114
rect 35 102 40 104
rect 60 103 64 113
rect 35 100 36 102
rect 38 100 40 102
rect 53 101 64 103
rect 35 98 50 100
rect 36 96 50 98
rect 53 99 54 101
rect 56 99 64 101
rect 53 97 64 99
rect 39 90 43 92
rect 39 88 40 90
rect 42 88 43 90
rect 39 82 43 88
rect 46 91 50 96
rect 84 93 88 113
rect 72 92 78 93
rect 46 90 61 91
rect 46 88 57 90
rect 59 88 61 90
rect 46 87 61 88
rect 72 90 74 92
rect 76 90 78 92
rect 72 82 78 90
rect 82 92 88 93
rect 82 90 84 92
rect 86 90 88 92
rect 82 89 88 90
rect 106 120 112 124
rect 128 123 168 124
rect 128 121 152 123
rect 154 121 168 123
rect 106 110 110 120
rect 116 119 120 121
rect 128 120 168 121
rect 116 117 117 119
rect 119 117 120 119
rect 116 116 120 117
rect 106 108 107 110
rect 109 108 110 110
rect 106 106 110 108
rect 113 112 120 116
rect 113 101 117 112
rect 156 107 160 112
rect 156 105 157 107
rect 159 105 160 107
rect 99 100 117 101
rect 99 98 101 100
rect 103 99 117 100
rect 103 98 128 99
rect 99 97 124 98
rect 113 96 124 97
rect 126 96 128 98
rect 113 95 128 96
rect 133 98 137 100
rect 133 96 134 98
rect 136 96 137 98
rect 133 91 137 96
rect 156 103 160 105
rect 164 109 168 120
rect 164 107 170 109
rect 164 105 167 107
rect 169 105 170 107
rect 164 103 170 105
rect 164 100 168 103
rect 148 96 168 100
rect 148 92 152 96
rect 112 90 134 91
rect 103 87 107 89
rect 112 88 114 90
rect 116 89 134 90
rect 136 89 137 91
rect 116 88 137 89
rect 142 91 152 92
rect 142 89 144 91
rect 146 89 152 91
rect 142 88 152 89
rect 197 124 221 128
rect 240 124 244 128
rect 195 120 201 124
rect 217 123 257 124
rect 217 121 241 123
rect 243 121 257 123
rect 195 110 199 120
rect 205 119 209 121
rect 217 120 257 121
rect 205 117 206 119
rect 208 117 209 119
rect 205 116 209 117
rect 195 108 196 110
rect 198 108 199 110
rect 195 106 199 108
rect 202 112 209 116
rect 202 101 206 112
rect 245 107 249 112
rect 245 105 246 107
rect 248 105 249 107
rect 188 100 206 101
rect 188 98 190 100
rect 192 99 206 100
rect 192 98 217 99
rect 188 97 213 98
rect 202 96 213 97
rect 215 96 217 98
rect 202 95 217 96
rect 222 98 226 100
rect 222 96 223 98
rect 225 96 226 98
rect 222 91 226 96
rect 245 103 249 105
rect 253 109 257 120
rect 283 124 287 128
rect 283 120 298 124
rect 253 107 259 109
rect 253 105 256 107
rect 258 105 259 107
rect 253 103 259 105
rect 253 100 257 103
rect 237 96 257 100
rect 237 92 241 96
rect 273 111 279 112
rect 294 107 298 120
rect 301 117 302 128
rect 324 130 330 138
rect 324 128 326 130
rect 328 128 330 130
rect 324 127 330 128
rect 358 130 364 138
rect 407 136 408 138
rect 410 136 411 138
rect 358 128 360 130
rect 362 128 364 130
rect 358 127 364 128
rect 294 105 295 107
rect 297 105 298 107
rect 294 99 298 105
rect 280 98 298 99
rect 280 96 282 98
rect 284 96 298 98
rect 280 95 298 96
rect 341 124 347 125
rect 330 122 343 124
rect 345 122 347 124
rect 330 120 347 122
rect 407 131 411 136
rect 407 129 408 131
rect 410 129 411 131
rect 201 90 223 91
rect 112 87 137 88
rect 192 87 196 89
rect 201 88 203 90
rect 205 89 223 90
rect 225 89 226 91
rect 205 88 226 89
rect 231 91 241 92
rect 231 89 233 91
rect 235 89 241 91
rect 231 88 241 89
rect 330 117 334 120
rect 321 113 334 117
rect 346 116 374 117
rect 321 99 325 113
rect 346 115 370 116
rect 346 113 347 115
rect 349 114 370 115
rect 372 114 374 116
rect 349 113 374 114
rect 346 101 350 113
rect 339 99 350 101
rect 321 97 322 99
rect 324 97 336 99
rect 321 95 336 97
rect 339 97 340 99
rect 342 97 350 99
rect 339 95 350 97
rect 201 87 226 88
rect 325 90 329 92
rect 325 88 326 90
rect 328 88 329 90
rect 103 85 104 87
rect 106 85 107 87
rect 192 85 193 87
rect 195 85 196 87
rect 270 85 276 86
rect 103 82 107 85
rect 159 84 165 85
rect 159 82 161 84
rect 163 82 165 84
rect 192 82 196 85
rect 248 84 254 85
rect 248 82 250 84
rect 252 82 254 84
rect 270 83 272 85
rect 274 83 276 85
rect 270 82 276 83
rect 289 85 295 86
rect 289 83 291 85
rect 293 83 295 85
rect 289 82 295 83
rect 325 82 329 88
rect 332 91 336 95
rect 370 91 374 113
rect 407 127 411 129
rect 425 131 431 139
rect 425 129 427 131
rect 429 129 431 131
rect 425 128 431 129
rect 459 131 465 139
rect 459 129 461 131
rect 463 129 465 131
rect 459 128 465 129
rect 489 131 495 139
rect 489 129 491 131
rect 493 129 495 131
rect 489 128 495 129
rect 523 131 529 139
rect 523 129 525 131
rect 527 129 529 131
rect 523 128 529 129
rect 553 131 559 139
rect 553 129 555 131
rect 557 129 559 131
rect 553 128 559 129
rect 587 131 593 139
rect 619 137 621 139
rect 623 137 625 139
rect 619 136 625 137
rect 587 129 589 131
rect 591 129 593 131
rect 587 128 593 129
rect 442 125 448 126
rect 442 123 444 125
rect 446 123 459 125
rect 442 121 459 123
rect 455 118 459 121
rect 415 117 443 118
rect 415 115 417 117
rect 419 116 443 117
rect 419 115 440 116
rect 415 114 440 115
rect 442 114 443 116
rect 332 90 347 91
rect 332 88 343 90
rect 345 88 347 90
rect 332 87 347 88
rect 358 90 364 91
rect 358 88 360 90
rect 362 88 364 90
rect 358 82 364 88
rect 368 90 374 91
rect 368 88 370 90
rect 372 88 374 90
rect 368 87 374 88
rect 385 97 389 99
rect 385 95 386 97
rect 388 95 389 97
rect 385 83 389 95
rect 406 97 411 99
rect 406 95 407 97
rect 409 95 411 97
rect 406 93 411 95
rect 407 83 411 93
rect 415 92 419 114
rect 439 102 443 114
rect 455 114 468 118
rect 439 100 450 102
rect 464 100 468 114
rect 439 98 447 100
rect 449 98 450 100
rect 439 96 450 98
rect 453 98 465 100
rect 467 98 468 100
rect 453 96 468 98
rect 453 92 457 96
rect 415 91 421 92
rect 415 89 417 91
rect 419 89 421 91
rect 415 88 421 89
rect 425 91 431 92
rect 425 89 427 91
rect 429 89 431 91
rect 425 83 431 89
rect 442 91 457 92
rect 442 89 444 91
rect 446 89 457 91
rect 442 88 457 89
rect 460 91 464 93
rect 460 89 461 91
rect 463 89 464 91
rect 460 83 464 89
rect 506 125 512 126
rect 495 123 508 125
rect 510 123 512 125
rect 495 121 512 123
rect 570 125 576 126
rect 559 123 572 125
rect 574 123 576 125
rect 559 121 576 123
rect 623 132 643 133
rect 623 130 639 132
rect 641 130 643 132
rect 623 129 643 130
rect 495 118 499 121
rect 486 114 499 118
rect 511 117 539 118
rect 486 100 490 114
rect 511 116 535 117
rect 511 114 512 116
rect 514 115 535 116
rect 537 115 539 117
rect 514 114 539 115
rect 511 102 515 114
rect 504 100 515 102
rect 486 98 487 100
rect 489 98 501 100
rect 486 96 501 98
rect 504 98 505 100
rect 507 98 515 100
rect 504 96 515 98
rect 490 91 494 93
rect 490 89 491 91
rect 493 89 494 91
rect 490 83 494 89
rect 497 92 501 96
rect 535 92 539 114
rect 497 91 512 92
rect 497 89 508 91
rect 510 89 512 91
rect 497 88 512 89
rect 523 91 529 92
rect 523 89 525 91
rect 527 89 529 91
rect 523 83 529 89
rect 533 91 539 92
rect 533 89 535 91
rect 537 89 539 91
rect 533 88 539 89
rect 559 118 563 121
rect 550 114 563 118
rect 575 117 603 118
rect 550 100 554 114
rect 575 116 599 117
rect 575 114 576 116
rect 578 115 599 116
rect 601 115 603 117
rect 578 114 603 115
rect 575 102 579 114
rect 568 100 579 102
rect 550 98 551 100
rect 553 98 565 100
rect 550 96 565 98
rect 568 98 569 100
rect 571 98 579 100
rect 568 96 579 98
rect 554 91 558 93
rect 554 89 555 91
rect 557 89 558 91
rect 554 83 558 89
rect 561 92 565 96
rect 599 92 603 114
rect 561 91 576 92
rect 561 89 572 91
rect 574 89 576 91
rect 561 88 576 89
rect 587 91 593 92
rect 587 89 589 91
rect 591 89 593 91
rect 587 83 593 89
rect 597 91 603 92
rect 597 89 599 91
rect 601 89 603 91
rect 597 88 603 89
rect 611 126 612 129
rect 623 125 627 129
rect 615 121 627 125
rect 615 109 619 121
rect 615 107 616 109
rect 618 107 619 109
rect 615 102 619 107
rect 615 98 632 102
rect 617 94 623 95
rect 617 92 619 94
rect 621 92 623 94
rect 617 83 623 92
rect 628 94 632 98
rect 652 113 653 119
rect 656 118 660 139
rect 679 121 683 139
rect 679 119 680 121
rect 682 119 683 121
rect 656 117 664 118
rect 656 115 660 117
rect 662 115 664 117
rect 656 114 664 115
rect 668 117 674 118
rect 679 117 683 119
rect 668 115 670 117
rect 672 115 674 117
rect 668 109 674 115
rect 655 108 674 109
rect 655 106 657 108
rect 659 106 674 108
rect 655 105 674 106
rect 628 92 629 94
rect 631 92 632 94
rect 628 90 632 92
rect 637 94 643 95
rect 637 92 639 94
rect 641 92 643 94
rect 637 83 643 92
rect 652 94 653 96
rect 664 92 668 105
rect 664 91 683 92
rect 664 89 679 91
rect 681 89 683 91
rect 664 88 683 89
rect 5 57 24 58
rect 5 55 7 57
rect 9 55 24 57
rect 5 54 24 55
rect 20 41 24 54
rect 35 50 36 52
rect 45 54 51 63
rect 45 52 47 54
rect 49 52 51 54
rect 45 51 51 52
rect 56 54 60 56
rect 56 52 57 54
rect 59 52 60 54
rect 14 40 33 41
rect 14 38 29 40
rect 31 38 33 40
rect 14 37 33 38
rect 14 31 20 37
rect 14 29 16 31
rect 18 29 20 31
rect 5 27 9 29
rect 14 28 20 29
rect 24 31 32 32
rect 24 29 26 31
rect 28 29 32 31
rect 24 28 32 29
rect 5 25 6 27
rect 8 25 9 27
rect 5 7 9 25
rect 28 7 32 28
rect 35 27 36 33
rect 56 48 60 52
rect 65 54 71 63
rect 65 52 67 54
rect 69 52 71 54
rect 65 51 71 52
rect 56 44 73 48
rect 69 39 73 44
rect 69 37 70 39
rect 72 37 73 39
rect 69 25 73 37
rect 61 21 73 25
rect 61 17 65 21
rect 76 17 77 20
rect 85 57 91 58
rect 85 55 87 57
rect 89 55 91 57
rect 85 54 91 55
rect 95 57 101 63
rect 95 55 97 57
rect 99 55 101 57
rect 95 54 101 55
rect 112 57 127 58
rect 112 55 114 57
rect 116 55 127 57
rect 112 54 127 55
rect 85 32 89 54
rect 123 50 127 54
rect 130 57 134 63
rect 130 55 131 57
rect 133 55 134 57
rect 130 53 134 55
rect 109 48 120 50
rect 109 46 117 48
rect 119 46 120 48
rect 123 48 138 50
rect 123 46 135 48
rect 137 46 138 48
rect 109 44 120 46
rect 109 32 113 44
rect 85 31 110 32
rect 85 29 87 31
rect 89 30 110 31
rect 112 30 113 32
rect 89 29 113 30
rect 134 32 138 46
rect 85 28 113 29
rect 125 28 138 32
rect 125 25 129 28
rect 149 57 155 58
rect 149 55 151 57
rect 153 55 155 57
rect 149 54 155 55
rect 159 57 165 63
rect 159 55 161 57
rect 163 55 165 57
rect 159 54 165 55
rect 176 57 191 58
rect 176 55 178 57
rect 180 55 191 57
rect 176 54 191 55
rect 149 32 153 54
rect 187 50 191 54
rect 194 57 198 63
rect 194 55 195 57
rect 197 55 198 57
rect 194 53 198 55
rect 173 48 184 50
rect 173 46 181 48
rect 183 46 184 48
rect 187 48 202 50
rect 187 46 199 48
rect 201 46 202 48
rect 173 44 184 46
rect 173 32 177 44
rect 149 31 174 32
rect 149 29 151 31
rect 153 30 174 31
rect 176 30 177 32
rect 153 29 177 30
rect 198 32 202 46
rect 149 28 177 29
rect 189 28 202 32
rect 189 25 193 28
rect 45 16 65 17
rect 45 14 47 16
rect 49 14 65 16
rect 45 13 65 14
rect 112 23 129 25
rect 112 21 114 23
rect 116 21 129 23
rect 112 20 118 21
rect 176 23 193 25
rect 176 21 178 23
rect 180 21 193 23
rect 176 20 182 21
rect 224 57 228 63
rect 224 55 225 57
rect 227 55 228 57
rect 224 53 228 55
rect 231 57 246 58
rect 231 55 242 57
rect 244 55 246 57
rect 231 54 246 55
rect 257 57 263 63
rect 257 55 259 57
rect 261 55 263 57
rect 257 54 263 55
rect 267 57 273 58
rect 267 55 269 57
rect 271 55 273 57
rect 267 54 273 55
rect 231 50 235 54
rect 220 48 235 50
rect 220 46 221 48
rect 223 46 235 48
rect 238 48 249 50
rect 238 46 239 48
rect 241 46 249 48
rect 220 32 224 46
rect 238 44 249 46
rect 220 28 233 32
rect 245 32 249 44
rect 269 32 273 54
rect 277 53 281 63
rect 277 51 282 53
rect 277 49 279 51
rect 281 49 282 51
rect 277 47 282 49
rect 299 51 303 63
rect 299 49 300 51
rect 302 49 303 51
rect 299 47 303 49
rect 314 58 320 59
rect 314 56 316 58
rect 318 56 320 58
rect 314 55 320 56
rect 324 58 330 64
rect 324 56 326 58
rect 328 56 330 58
rect 324 55 330 56
rect 341 58 356 59
rect 341 56 343 58
rect 345 56 356 58
rect 341 55 356 56
rect 245 30 246 32
rect 248 31 273 32
rect 248 30 269 31
rect 245 29 269 30
rect 271 29 273 31
rect 245 28 273 29
rect 229 25 233 28
rect 229 23 246 25
rect 229 21 242 23
rect 244 21 246 23
rect 240 20 246 21
rect 95 17 101 18
rect 95 15 97 17
rect 99 15 101 17
rect 63 9 69 10
rect 63 7 65 9
rect 67 7 69 9
rect 95 7 101 15
rect 129 17 135 18
rect 129 15 131 17
rect 133 15 135 17
rect 129 7 135 15
rect 159 17 165 18
rect 159 15 161 17
rect 163 15 165 17
rect 159 7 165 15
rect 193 17 199 18
rect 193 15 195 17
rect 197 15 199 17
rect 193 7 199 15
rect 223 17 229 18
rect 223 15 225 17
rect 227 15 229 17
rect 223 7 229 15
rect 257 17 263 18
rect 257 15 259 17
rect 261 15 263 17
rect 257 7 263 15
rect 277 17 281 19
rect 314 33 318 55
rect 352 51 356 55
rect 359 58 363 64
rect 393 63 399 64
rect 393 61 395 63
rect 397 61 399 63
rect 393 60 399 61
rect 412 63 418 64
rect 412 61 414 63
rect 416 61 418 63
rect 434 62 436 64
rect 438 62 440 64
rect 434 61 440 62
rect 492 61 496 64
rect 523 62 525 64
rect 527 62 529 64
rect 523 61 529 62
rect 581 61 585 64
rect 412 60 418 61
rect 492 59 493 61
rect 495 59 496 61
rect 581 59 582 61
rect 584 59 585 61
rect 359 56 360 58
rect 362 56 363 58
rect 359 54 363 56
rect 462 58 487 59
rect 338 49 349 51
rect 338 47 346 49
rect 348 47 349 49
rect 352 49 367 51
rect 352 47 364 49
rect 366 47 367 49
rect 338 45 349 47
rect 338 33 342 45
rect 314 32 339 33
rect 314 30 316 32
rect 318 31 339 32
rect 341 31 342 33
rect 318 30 342 31
rect 363 33 367 47
rect 314 29 342 30
rect 354 29 367 33
rect 354 26 358 29
rect 447 57 457 58
rect 447 55 453 57
rect 455 55 457 57
rect 447 54 457 55
rect 462 57 483 58
rect 462 55 463 57
rect 465 56 483 57
rect 485 56 487 58
rect 492 57 496 59
rect 551 58 576 59
rect 465 55 487 56
rect 277 15 278 17
rect 280 15 281 17
rect 277 10 281 15
rect 341 24 358 26
rect 341 22 343 24
rect 345 22 358 24
rect 341 21 347 22
rect 390 50 408 51
rect 390 48 404 50
rect 406 48 408 50
rect 390 47 408 48
rect 390 41 394 47
rect 390 39 391 41
rect 393 39 394 41
rect 324 18 330 19
rect 324 16 326 18
rect 328 16 330 18
rect 277 8 278 10
rect 280 8 281 10
rect 324 8 330 16
rect 358 18 364 19
rect 358 16 360 18
rect 362 16 364 18
rect 358 8 364 16
rect 386 18 387 29
rect 390 26 394 39
rect 409 34 415 35
rect 447 50 451 54
rect 431 46 451 50
rect 431 43 435 46
rect 429 41 435 43
rect 429 39 430 41
rect 432 39 435 41
rect 429 37 435 39
rect 390 22 405 26
rect 401 18 405 22
rect 431 26 435 37
rect 439 41 443 43
rect 462 50 466 55
rect 462 48 463 50
rect 465 48 466 50
rect 462 46 466 48
rect 471 50 486 51
rect 471 48 473 50
rect 475 49 486 50
rect 475 48 500 49
rect 471 47 496 48
rect 482 46 496 47
rect 498 46 500 48
rect 482 45 500 46
rect 439 39 440 41
rect 442 39 443 41
rect 439 34 443 39
rect 482 34 486 45
rect 479 30 486 34
rect 489 38 493 40
rect 489 36 490 38
rect 492 36 493 38
rect 479 29 483 30
rect 479 27 480 29
rect 482 27 483 29
rect 431 25 471 26
rect 479 25 483 27
rect 489 26 493 36
rect 431 23 445 25
rect 447 23 471 25
rect 431 22 471 23
rect 487 22 493 26
rect 444 18 448 22
rect 467 18 491 22
rect 536 57 546 58
rect 536 55 542 57
rect 544 55 546 57
rect 536 54 546 55
rect 551 57 572 58
rect 551 55 552 57
rect 554 56 572 57
rect 574 56 576 58
rect 581 57 585 59
rect 554 55 576 56
rect 536 50 540 54
rect 520 46 540 50
rect 520 43 524 46
rect 518 41 524 43
rect 518 39 519 41
rect 521 39 524 41
rect 518 37 524 39
rect 520 26 524 37
rect 528 41 532 43
rect 551 50 555 55
rect 551 48 552 50
rect 554 48 555 50
rect 551 46 555 48
rect 560 50 575 51
rect 560 48 562 50
rect 564 49 575 50
rect 564 48 589 49
rect 560 47 585 48
rect 571 46 585 47
rect 587 46 589 48
rect 571 45 589 46
rect 528 39 529 41
rect 531 39 532 41
rect 528 34 532 39
rect 571 34 575 45
rect 568 30 575 34
rect 578 38 582 40
rect 578 36 579 38
rect 581 36 582 38
rect 568 29 572 30
rect 568 27 569 29
rect 571 27 572 29
rect 520 25 560 26
rect 568 25 572 27
rect 578 26 582 36
rect 520 23 534 25
rect 536 23 560 25
rect 520 22 560 23
rect 576 22 582 26
rect 600 56 606 57
rect 600 54 602 56
rect 604 54 606 56
rect 600 53 606 54
rect 610 56 616 64
rect 610 54 612 56
rect 614 54 616 56
rect 627 58 642 59
rect 627 56 629 58
rect 631 56 642 58
rect 627 55 642 56
rect 610 53 616 54
rect 600 33 604 53
rect 638 50 642 55
rect 645 58 649 64
rect 645 56 646 58
rect 648 56 649 58
rect 645 54 649 56
rect 624 47 635 49
rect 624 45 632 47
rect 634 45 635 47
rect 638 48 652 50
rect 638 46 653 48
rect 624 43 635 45
rect 648 44 650 46
rect 652 44 653 46
rect 624 33 628 43
rect 648 42 653 44
rect 600 32 628 33
rect 600 30 602 32
rect 604 31 628 32
rect 604 30 625 31
rect 600 29 625 30
rect 627 29 628 31
rect 644 32 645 38
rect 624 27 628 29
rect 533 18 537 22
rect 556 18 580 22
rect 401 17 418 18
rect 401 15 414 17
rect 416 15 418 17
rect 401 14 418 15
rect 433 17 439 18
rect 433 15 435 17
rect 437 15 439 17
rect 393 10 399 11
rect 393 8 395 10
rect 397 8 399 10
rect 433 10 439 15
rect 444 16 445 18
rect 447 16 448 18
rect 444 14 448 16
rect 455 17 461 18
rect 455 15 457 17
rect 459 15 461 17
rect 433 8 435 10
rect 437 8 439 10
rect 455 10 461 15
rect 522 17 528 18
rect 522 15 524 17
rect 526 15 528 17
rect 455 8 457 10
rect 459 8 461 10
rect 490 10 496 11
rect 490 8 492 10
rect 494 8 496 10
rect 522 10 528 15
rect 533 16 534 18
rect 536 16 537 18
rect 533 14 537 16
rect 544 17 550 18
rect 544 15 546 17
rect 548 15 550 17
rect 522 8 524 10
rect 526 8 528 10
rect 544 10 550 15
rect 648 25 652 42
rect 636 21 652 25
rect 627 20 640 21
rect 627 18 629 20
rect 631 18 640 20
rect 679 53 683 64
rect 668 46 669 52
rect 679 51 680 53
rect 682 51 683 53
rect 679 49 683 51
rect 668 27 669 34
rect 627 17 640 18
rect 675 17 681 18
rect 675 15 677 17
rect 679 15 681 17
rect 544 8 546 10
rect 548 8 550 10
rect 579 10 585 11
rect 579 8 581 10
rect 583 8 585 10
rect 611 10 615 12
rect 611 8 612 10
rect 614 8 615 10
rect 644 10 650 11
rect 644 8 646 10
rect 648 8 650 10
rect 675 8 681 15
<< via1 >>
rect 6 252 8 254
rect 21 247 23 249
rect 29 252 31 254
rect 49 260 51 262
rect 69 244 71 246
rect 152 260 154 262
rect 93 240 95 242
rect 141 243 143 245
rect 174 243 176 245
rect 182 260 184 262
rect 214 252 216 254
rect 370 276 372 278
rect 303 254 305 256
rect 271 243 273 245
rect 339 254 341 256
rect 360 243 362 245
rect 416 276 418 278
rect 536 275 538 277
rect 600 276 602 278
rect 401 269 403 271
rect 385 257 387 259
rect 409 261 411 263
rect 429 245 431 247
rect 452 254 454 256
rect 472 254 474 256
rect 500 254 502 256
rect 524 245 526 247
rect 544 245 546 247
rect 569 257 571 259
rect 592 244 594 246
rect 608 257 610 259
rect 632 270 634 272
rect 640 253 642 255
rect 665 270 667 272
rect 681 253 683 255
rect 649 244 651 246
rect 37 194 39 196
rect 5 185 7 187
rect 21 168 23 170
rect 46 185 48 187
rect 54 168 56 170
rect 78 181 80 183
rect 94 194 96 196
rect 117 181 119 183
rect 142 193 144 195
rect 162 193 164 195
rect 186 184 188 186
rect 214 184 216 186
rect 234 184 236 186
rect 257 193 259 195
rect 277 177 279 179
rect 301 181 303 183
rect 285 169 287 171
rect 86 162 88 164
rect 150 163 152 165
rect 270 162 272 164
rect 326 195 328 197
rect 347 184 349 186
rect 371 176 373 178
rect 415 195 417 197
rect 383 184 385 186
rect 316 162 318 164
rect 472 186 474 188
rect 504 178 506 180
rect 512 195 514 197
rect 545 195 547 197
rect 593 198 595 200
rect 534 178 536 180
rect 617 194 619 196
rect 637 178 639 180
rect 602 169 604 171
rect 657 186 659 188
rect 665 191 667 193
rect 680 186 682 188
rect 6 105 8 107
rect 21 100 23 102
rect 29 105 31 107
rect 49 113 51 115
rect 69 97 71 99
rect 152 113 154 115
rect 93 93 95 95
rect 141 96 143 98
rect 174 96 176 98
rect 182 113 184 115
rect 214 105 216 107
rect 370 129 372 131
rect 303 107 305 109
rect 271 96 273 98
rect 339 107 341 109
rect 360 96 362 98
rect 416 129 418 131
rect 536 128 538 130
rect 600 129 602 131
rect 401 122 403 124
rect 385 110 387 112
rect 409 114 411 116
rect 429 98 431 100
rect 452 107 454 109
rect 472 107 474 109
rect 500 107 502 109
rect 524 98 526 100
rect 544 98 546 100
rect 569 110 571 112
rect 592 97 594 99
rect 608 110 610 112
rect 632 123 634 125
rect 640 106 642 108
rect 665 123 667 125
rect 681 106 683 108
rect 649 97 651 99
rect 37 47 39 49
rect 5 38 7 40
rect 21 21 23 23
rect 46 38 48 40
rect 54 21 56 23
rect 78 34 80 36
rect 94 47 96 49
rect 117 34 119 36
rect 142 46 144 48
rect 162 46 164 48
rect 186 37 188 39
rect 214 37 216 39
rect 234 37 236 39
rect 257 46 259 48
rect 277 30 279 32
rect 301 34 303 36
rect 285 22 287 24
rect 86 15 88 17
rect 150 16 152 18
rect 270 15 272 17
rect 326 48 328 50
rect 347 37 349 39
rect 415 48 417 50
rect 383 37 385 39
rect 316 15 318 17
rect 472 39 474 41
rect 504 31 506 33
rect 512 48 514 50
rect 545 48 547 50
rect 593 51 595 53
rect 534 31 536 33
rect 617 47 619 49
rect 637 31 639 33
rect 657 39 659 41
rect 602 16 604 18
rect 665 44 667 46
rect 680 39 682 41
<< via2 >>
rect 178 243 180 245
rect 472 276 474 278
rect 535 268 537 270
rect 623 261 625 263
rect 63 177 65 179
rect 545 202 547 204
rect 508 195 510 197
rect 377 176 379 178
rect 602 161 604 163
rect 178 96 180 98
rect 471 129 473 131
rect 535 121 537 123
rect 623 114 625 116
rect 424 98 426 100
rect 63 30 65 32
rect 508 48 510 50
rect 602 22 604 24
rect 602 13 604 15
<< via3 >>
rect 476 276 478 278
rect 536 278 538 280
rect 598 161 600 163
rect 476 129 478 131
rect 536 131 538 133
rect 606 23 608 25
<< labels >>
rlabel alu1 510 68 510 68 5 Vss
rlabel alu1 510 4 510 4 5 Vdd
rlabel alu1 344 4 344 4 2 vdd
rlabel alu1 344 68 344 68 2 vss
rlabel alu1 445 79 445 79 4 vss
rlabel alu1 445 143 445 143 4 vdd
rlabel alu1 509 79 509 79 6 vss
rlabel alu1 509 143 509 143 6 vdd
rlabel alu1 573 143 573 143 6 vdd
rlabel alu1 573 79 573 79 6 vss
rlabel alu1 666 143 666 143 6 vdd
rlabel alu1 625 79 625 79 6 vss
rlabel alu1 625 143 625 143 6 vdd
rlabel space 605 78 645 146 1 or
rlabel space 647 78 687 146 1 and
rlabel space 408 78 605 146 1 4x1_mux
rlabel alu1 666 79 666 79 6 vss
rlabel space 377 0 688 76 1 fafs
rlabel space 312 0 376 76 1 shift_mux
rlabel alu1 398 78 398 78 6 vss
rlabel alu1 398 142 398 142 6 vdd
rlabel ab 383 77 412 146 1 decoder
rlabel alu1 536 133 536 133 1 s1
rlabel alu2 475 130 475 130 1 s0
rlabel alu1 178 78 178 78 1 Vss
rlabel alu1 30 120 30 120 1 b_test
rlabel alu1 75 98 75 98 1 Bn
rlabel alu1 86 132 86 132 1 Binv
rlabel alu1 94 109 94 109 1 Sum
rlabel via1 50 114 50 114 1 B
rlabel alu1 231 96 231 96 1 A
rlabel alu1 178 142 178 142 1 Vdd
rlabel alu1 142 98 142 98 1 Cin
rlabel alu1 316 110 316 110 5 COUT
rlabel alu1 344 142 344 142 6 vdd
rlabel alu1 344 78 344 78 6 vss
rlabel alu1 304 111 304 111 5 fafs_cout
rlabel via1 361 97 361 97 5 in1
rlabel alu2 336 109 336 109 5 in2
rlabel alu1 231 39 231 39 8 a0
rlabel alu1 243 67 243 67 8 vss
rlabel alu1 255 43 255 43 8 a1
rlabel alu1 243 3 243 3 8 vdd
rlabel via1 215 39 215 39 5 y0
rlabel alu1 179 67 179 67 2 vss
rlabel alu1 179 3 179 3 2 vdd
rlabel alu2 166 47 166 47 5 k1
rlabel alu1 143 38 144 40 5 y1
rlabel alu1 99 47 99 47 5 a3
rlabel alu1 115 3 115 3 2 vdd
rlabel alu1 115 67 115 67 2 vss
rlabel alu1 263 47 263 47 8 a1
rlabel alu1 22 19 22 19 2 a
rlabel alu1 14 47 14 47 2 b
rlabel alu1 14 15 14 15 2 a
rlabel alu1 22 3 22 3 2 vdd
rlabel alu1 207 42 207 42 5 out
rlabel alu1 63 67 63 67 2 vss
rlabel alu1 63 31 63 31 2 a
rlabel alu1 63 3 63 3 2 vdd
rlabel alu1 55 39 55 39 2 b
rlabel alu1 55 23 55 23 2 a
rlabel space 43 0 83 68 5 or
rlabel space 1 0 41 68 5 and
rlabel alu1 47 35 47 35 2 b
rlabel alu4 38 48 38 48 5 z3
rlabel via1 79 35 79 35 5 z2
rlabel space 83 0 280 68 5 4x1_mux
rlabel via1 188 37 188 37 5 k0
rlabel alu1 6 43 6 43 2 b
rlabel alu1 22 67 22 67 2 vss
rlabel space 0 70 311 146 5 fafs
rlabel space 312 70 376 146 5 shift_mux
rlabel alu1 372 130 372 130 7 fafs_en
rlabel alu1 302 28 302 28 2 z
rlabel alu1 294 48 294 48 2 z
rlabel alu1 290 68 290 68 2 vss
rlabel alu1 290 4 290 4 2 vdd
rlabel alu1 282 40 282 40 5 l1
rlabel alu1 291 28 291 28 5 l0
rlabel ab 276 0 305 69 5 decoder
rlabel alu1 124 38 124 38 5 or_out
rlabel alu1 152 13 152 13 5 s1
rlabel alu2 213 16 213 16 5 s0
rlabel alu1 178 225 178 225 1 Vss
rlabel alu1 30 267 30 267 1 b_test
rlabel alu1 75 245 75 245 1 Bn
rlabel alu1 86 279 86 279 1 Binv
rlabel alu1 94 256 94 256 1 Sum
rlabel via1 50 261 50 261 1 B
rlabel alu1 231 243 231 243 1 A
rlabel alu1 178 289 178 289 1 Vdd
rlabel alu1 142 245 142 245 1 Cin
rlabel alu1 316 257 316 257 5 COUT
rlabel alu1 344 289 344 289 6 vdd
rlabel alu1 344 225 344 225 6 vss
rlabel alu1 304 258 304 258 5 fafs_cout
rlabel via1 361 244 361 244 5 in1
rlabel alu2 336 256 336 256 5 in2
rlabel alu1 231 186 231 186 8 a0
rlabel alu1 243 214 243 214 8 vss
rlabel alu1 255 190 255 190 8 a1
rlabel alu1 243 150 243 150 8 vdd
rlabel via1 215 186 215 186 5 y0
rlabel alu1 179 214 179 214 2 vss
rlabel alu1 179 150 179 150 2 vdd
rlabel alu2 166 194 166 194 5 k1
rlabel alu1 143 185 144 187 5 y1
rlabel alu1 99 194 99 194 5 a3
rlabel alu1 115 150 115 150 2 vdd
rlabel alu1 115 214 115 214 2 vss
rlabel alu1 263 194 263 194 8 a1
rlabel alu1 22 166 22 166 2 a
rlabel alu1 14 194 14 194 2 b
rlabel alu1 14 162 14 162 2 a
rlabel alu1 22 150 22 150 2 vdd
rlabel alu1 207 189 207 189 5 out
rlabel alu1 63 214 63 214 2 vss
rlabel alu1 63 178 63 178 2 a
rlabel alu1 63 150 63 150 2 vdd
rlabel alu1 55 186 55 186 2 b
rlabel alu1 55 170 55 170 2 a
rlabel space 43 147 83 215 5 or
rlabel space 1 147 41 215 5 and
rlabel alu1 47 182 47 182 2 b
rlabel alu4 38 195 38 195 5 z3
rlabel via1 79 182 79 182 5 z2
rlabel space 83 147 280 215 5 4x1_mux
rlabel via1 188 184 188 184 5 k0
rlabel alu1 6 190 6 190 2 b
rlabel alu1 22 214 22 214 2 vss
rlabel space 0 217 311 293 5 fafs
rlabel space 312 217 376 293 5 shift_mux
rlabel alu1 372 277 372 277 7 fafs_en
rlabel alu1 302 175 302 175 2 z
rlabel alu1 294 195 294 195 2 z
rlabel alu1 290 215 290 215 2 vss
rlabel alu1 290 151 290 151 2 vdd
rlabel alu1 282 187 282 187 5 l1
rlabel alu1 291 175 291 175 5 l0
rlabel ab 276 147 305 216 5 decoder
rlabel alu1 124 185 124 185 5 or_out
rlabel alu1 152 160 152 160 5 s1
rlabel alu2 213 163 213 163 5 s0
rlabel alu1 510 215 510 215 5 Vss
rlabel alu1 510 151 510 151 5 Vdd
rlabel alu1 344 151 344 151 2 vdd
rlabel alu1 344 215 344 215 2 vss
rlabel alu1 445 226 445 226 4 vss
rlabel alu1 445 290 445 290 4 vdd
rlabel alu1 509 226 509 226 6 vss
rlabel alu1 509 290 509 290 6 vdd
rlabel alu1 573 290 573 290 6 vdd
rlabel alu1 573 226 573 226 6 vss
rlabel alu1 666 290 666 290 6 vdd
rlabel alu1 625 226 625 226 6 vss
rlabel alu1 625 290 625 290 6 vdd
rlabel space 605 225 645 293 1 or
rlabel space 647 225 687 293 1 and
rlabel space 408 225 605 293 1 4x1_mux
rlabel alu1 666 226 666 226 6 vss
rlabel space 377 147 688 223 1 fafs
rlabel space 312 147 376 223 1 shift_mux
rlabel alu1 316 163 316 163 3 fafs_en
rlabel alu1 398 225 398 225 6 vss
rlabel alu1 398 289 398 289 6 vdd
rlabel ab 383 224 412 293 1 decoder
rlabel alu1 536 280 536 280 1 s1
rlabel alu2 475 277 475 277 1 s0
rlabel via1 638 180 638 180 1 B0
rlabel alu1 372 182 372 182 1 COUT0
rlabel alu2 458 48 458 48 1 A1
rlabel alu1 372 34 372 34 1 COUT1
rlabel alu2 546 46 546 46 1 CIN1
rlabel via1 638 31 638 31 1 B1
rlabel alu1 602 15 602 15 1 BINV
rlabel alu1 481 104 481 104 1 OUT1
rlabel alu1 481 251 481 251 1 OUT0
rlabel alu1 593 47 593 47 1 SUM
rlabel alu1 594 192 594 192 1 SUM0
rlabel via2 602 161 602 161 1 B_INV
rlabel alu3 546 200 546 200 1 CIN0
rlabel alu1 691 249 691 249 1 B0
rlabel alu1 689 279 689 279 1 A0
<< end >>
